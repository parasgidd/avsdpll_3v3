magic
tech scmos
timestamp 1627569390
<< nwell >>
rect 550 550 579 593
rect 632 550 687 593
rect 760 550 814 593
<< ntransistor >>
rect 561 489 563 492
rect 653 487 655 493
rect 663 487 665 493
rect 775 484 777 493
rect 786 484 788 493
rect 797 484 799 493
<< ptransistor >>
rect 561 556 563 567
rect 653 556 655 567
rect 663 556 665 567
rect 775 556 777 567
rect 786 556 788 567
rect 797 556 799 567
<< ndiffusion >>
rect 560 489 561 492
rect 563 489 564 492
rect 651 487 653 493
rect 655 487 663 493
rect 665 487 667 493
rect 773 484 775 493
rect 777 484 786 493
rect 788 484 797 493
rect 799 484 801 493
<< pdiffusion >>
rect 560 556 561 567
rect 563 556 564 567
rect 651 556 653 567
rect 655 556 657 567
rect 661 556 663 567
rect 665 556 667 567
rect 773 556 775 567
rect 777 556 780 567
rect 784 556 786 567
rect 788 556 791 567
rect 795 556 797 567
rect 799 556 801 567
<< ndcontact >>
rect 556 488 560 493
rect 564 488 568 493
rect 647 487 651 493
rect 667 487 671 493
rect 769 484 773 493
rect 801 484 805 493
<< pdcontact >>
rect 556 556 560 567
rect 564 556 568 567
rect 647 556 651 567
rect 657 556 661 567
rect 667 556 671 567
rect 769 556 773 567
rect 780 556 784 567
rect 791 556 795 567
rect 801 556 805 567
<< psubstratepcontact >>
rect 559 472 563 476
rect 567 472 571 476
rect 642 472 646 476
rect 650 472 654 476
rect 658 472 662 476
rect 666 472 670 476
rect 674 472 678 476
rect 768 472 772 476
rect 776 472 780 476
rect 784 472 788 476
rect 792 472 796 476
rect 800 472 804 476
<< nsubstratencontact >>
rect 553 582 557 586
rect 561 582 565 586
rect 569 582 573 586
rect 638 582 642 586
rect 646 582 650 586
rect 655 582 659 586
rect 663 582 667 586
rect 671 582 675 586
rect 769 582 773 586
rect 777 582 781 586
rect 787 582 791 586
rect 795 582 799 586
rect 553 574 557 578
rect 561 574 565 578
rect 569 574 573 578
rect 638 574 642 578
rect 646 574 650 578
rect 655 574 659 578
rect 663 574 667 578
rect 671 574 675 578
rect 769 574 773 578
rect 777 574 781 578
rect 787 574 791 578
rect 795 574 799 578
<< polysilicon >>
rect 561 567 563 569
rect 653 567 655 569
rect 663 567 665 569
rect 775 567 777 569
rect 786 567 788 569
rect 797 567 799 569
rect 561 492 563 556
rect 653 493 655 556
rect 663 511 665 556
rect 775 537 777 556
rect 663 493 665 506
rect 775 493 777 532
rect 786 526 788 556
rect 797 531 799 556
rect 787 521 788 526
rect 786 493 788 521
rect 797 493 799 526
rect 561 487 563 489
rect 653 485 655 487
rect 663 485 665 487
rect 775 482 777 484
rect 786 482 788 484
rect 797 482 799 484
<< polycontact >>
rect 556 520 561 525
rect 648 496 653 501
rect 774 532 779 537
rect 660 506 665 511
rect 795 526 799 531
rect 782 521 787 526
<< metal1 >>
rect 550 586 579 587
rect 550 582 553 586
rect 557 582 561 586
rect 565 582 569 586
rect 573 582 579 586
rect 550 578 579 582
rect 550 574 553 578
rect 557 574 561 578
rect 565 574 569 578
rect 573 574 579 578
rect 550 573 579 574
rect 632 586 687 587
rect 632 582 638 586
rect 642 582 646 586
rect 650 582 655 586
rect 659 582 663 586
rect 667 582 671 586
rect 675 582 687 586
rect 632 578 687 582
rect 632 574 638 578
rect 642 574 646 578
rect 650 574 655 578
rect 659 574 663 578
rect 667 574 671 578
rect 675 574 687 578
rect 632 573 687 574
rect 760 586 814 587
rect 760 582 769 586
rect 773 582 777 586
rect 781 582 787 586
rect 791 582 795 586
rect 799 582 814 586
rect 760 578 814 582
rect 760 574 769 578
rect 773 574 777 578
rect 781 574 787 578
rect 791 574 795 578
rect 799 574 814 578
rect 760 573 814 574
rect 556 567 559 573
rect 647 567 650 573
rect 668 567 671 573
rect 769 567 772 573
rect 791 567 794 573
rect 565 534 568 556
rect 565 531 573 534
rect 553 521 556 524
rect 565 493 568 531
rect 657 520 660 556
rect 780 544 783 556
rect 802 544 805 556
rect 780 541 812 544
rect 760 533 774 536
rect 760 522 782 525
rect 657 517 678 520
rect 638 507 660 510
rect 638 497 648 500
rect 668 493 671 517
rect 802 493 805 541
rect 556 479 559 488
rect 647 479 650 487
rect 769 479 772 484
rect 550 476 579 479
rect 550 472 559 476
rect 563 472 567 476
rect 571 472 579 476
rect 550 469 579 472
rect 632 476 687 479
rect 632 472 642 476
rect 646 472 650 476
rect 654 472 658 476
rect 662 472 666 476
rect 670 472 674 476
rect 678 472 687 476
rect 632 469 687 472
rect 760 476 814 479
rect 760 472 768 476
rect 772 472 776 476
rect 780 472 784 476
rect 788 472 792 476
rect 796 472 800 476
rect 804 472 814 476
rect 760 469 814 472
<< m2contact >>
rect 795 526 799 531
<< metal2 >>
rect 760 528 795 531
<< end >>
