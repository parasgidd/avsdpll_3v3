magic
tech scmos
timestamp 1598358295
<< nwell >>
rect -4 -27 158 -2
<< ntransistor >>
rect 10 50 12 53
rect 29 50 31 53
rect 49 50 51 53
rect 61 50 63 53
rect 79 50 81 53
rect 95 50 97 53
rect 109 50 111 53
rect 122 50 124 53
rect 143 50 145 53
<< ptransistor >>
rect 10 -16 12 -8
rect 29 -16 31 -8
rect 49 -16 51 -8
rect 61 -16 63 -8
rect 79 -16 81 -8
rect 95 -16 97 -8
rect 109 -16 111 -8
rect 122 -16 124 -8
rect 143 -16 145 -8
<< ndiffusion >>
rect 7 50 10 53
rect 12 50 13 53
rect 27 50 29 53
rect 31 50 32 53
rect 46 50 49 53
rect 51 50 54 53
rect 59 50 61 53
rect 63 50 64 53
rect 78 50 79 53
rect 81 50 86 53
rect 91 50 95 53
rect 97 50 101 53
rect 106 50 109 53
rect 111 50 114 53
rect 119 50 122 53
rect 124 50 127 53
rect 141 50 143 53
rect 145 50 146 53
<< pdiffusion >>
rect 7 -16 10 -8
rect 12 -16 13 -8
rect 27 -16 29 -8
rect 31 -16 32 -8
rect 46 -16 49 -8
rect 51 -16 54 -8
rect 59 -16 61 -8
rect 63 -16 64 -8
rect 78 -16 79 -8
rect 81 -16 86 -8
rect 91 -16 95 -8
rect 97 -16 101 -8
rect 106 -16 109 -8
rect 111 -16 114 -8
rect 119 -16 122 -8
rect 124 -16 127 -8
rect 141 -16 143 -8
rect 145 -16 146 -8
<< ndcontact >>
rect 2 49 7 54
rect 13 49 18 54
rect 22 49 27 54
rect 32 49 37 54
rect 41 49 46 54
rect 54 49 59 54
rect 64 49 69 54
rect 73 49 78 54
rect 86 49 91 54
rect 101 49 106 54
rect 114 49 119 54
rect 127 49 132 54
rect 136 49 141 54
rect 146 49 151 54
<< pdcontact >>
rect 2 -16 7 -8
rect 13 -16 18 -8
rect 22 -16 27 -8
rect 32 -16 37 -8
rect 41 -16 46 -8
rect 54 -16 59 -8
rect 64 -16 69 -8
rect 73 -16 78 -8
rect 86 -16 91 -8
rect 101 -16 106 -8
rect 114 -16 119 -8
rect 127 -16 132 -8
rect 136 -16 141 -8
rect 146 -16 151 -8
<< psubstratepcontact >>
rect -2 80 3 85
rect 7 80 12 85
rect 16 80 21 85
rect 25 80 30 85
rect 35 80 40 85
rect 44 80 49 85
rect 54 80 59 85
rect 63 80 68 85
rect 74 80 79 85
rect 84 80 89 85
rect 93 80 98 85
rect 102 80 107 85
rect 111 80 116 85
rect 120 80 125 85
rect 129 80 134 85
rect 138 80 143 85
rect 147 80 152 85
rect -2 71 3 76
rect 7 71 12 76
rect 16 71 21 76
rect 25 71 30 76
rect 35 71 40 76
rect 44 71 49 76
rect 54 71 59 76
rect 63 71 68 76
rect 74 71 79 76
rect 84 71 89 76
rect 93 71 98 76
rect 102 71 107 76
rect 111 71 116 76
rect 120 71 125 76
rect 129 71 134 76
rect 138 71 143 76
rect 147 71 152 76
<< nsubstratencontact >>
rect -2 -42 3 -37
rect 7 -42 12 -37
rect 17 -42 22 -37
rect 26 -42 31 -37
rect 35 -42 40 -37
rect 44 -42 49 -37
rect 53 -42 58 -37
rect 62 -42 67 -37
rect 72 -42 77 -37
rect 81 -42 86 -37
rect 91 -42 96 -37
rect 101 -42 106 -37
rect 111 -42 116 -37
rect 120 -42 125 -37
rect 130 -42 135 -37
rect 139 -42 144 -37
rect 148 -42 153 -37
rect -2 -51 3 -46
rect 7 -51 12 -46
rect 17 -51 22 -46
rect 26 -51 31 -46
rect 35 -51 40 -46
rect 44 -51 49 -46
rect 53 -51 58 -46
rect 62 -51 67 -46
rect 72 -51 77 -46
rect 81 -51 86 -46
rect 91 -51 96 -46
rect 101 -51 106 -46
rect 111 -51 116 -46
rect 120 -51 125 -46
rect 130 -51 135 -46
rect 139 -51 144 -46
rect 148 -51 153 -46
<< polysilicon >>
rect 10 53 12 55
rect 10 7 12 50
rect 29 53 31 55
rect 29 17 31 50
rect 49 53 51 55
rect 49 32 51 50
rect 61 53 63 55
rect 10 -8 12 2
rect 29 -8 31 12
rect 61 10 63 50
rect 79 53 81 55
rect 79 48 81 50
rect 95 53 97 55
rect 95 48 97 50
rect 109 53 111 55
rect 79 46 97 48
rect 109 33 111 50
rect 122 53 124 55
rect 122 24 124 50
rect 143 53 145 55
rect 143 32 145 50
rect 49 -8 51 -2
rect 61 -8 63 5
rect 79 -6 94 -4
rect 79 -8 81 -6
rect 95 -8 97 -6
rect 109 -8 111 -2
rect 122 -8 124 19
rect 143 -8 145 27
rect 10 -18 12 -16
rect 29 -18 31 -16
rect 49 -18 51 -16
rect 61 -18 63 -16
rect 79 -18 81 -16
rect 95 -18 97 -16
rect 109 -18 111 -16
rect 122 -18 124 -16
rect 143 -18 145 -16
<< polycontact >>
rect 48 27 52 32
rect 29 12 33 17
rect 10 2 14 7
rect 80 41 84 46
rect 108 28 112 33
rect 143 27 147 32
rect 122 19 126 24
rect 61 5 65 10
rect 48 -2 52 3
rect 94 -6 98 -1
rect 108 -2 112 3
<< metal1 >>
rect -4 85 157 89
rect -4 80 -2 85
rect 3 80 7 85
rect 12 80 16 85
rect 21 80 25 85
rect 30 80 35 85
rect 40 80 44 85
rect 49 80 54 85
rect 59 80 63 85
rect 68 80 74 85
rect 79 80 84 85
rect 89 80 93 85
rect 98 80 102 85
rect 107 80 111 85
rect 116 80 120 85
rect 125 80 129 85
rect 134 80 138 85
rect 143 80 147 85
rect 152 80 157 85
rect -4 76 157 80
rect -4 71 -2 76
rect 3 71 7 76
rect 12 71 16 76
rect 21 71 25 76
rect 30 71 35 76
rect 40 71 44 76
rect 49 71 54 76
rect 59 71 63 76
rect 68 71 74 76
rect 79 71 84 76
rect 89 71 93 76
rect 98 71 102 76
rect 107 71 111 76
rect 116 71 120 76
rect 125 71 129 76
rect 134 71 138 76
rect 143 71 147 76
rect 152 71 157 76
rect -4 69 157 71
rect 14 54 17 69
rect 33 54 36 69
rect 65 54 68 69
rect 128 54 131 69
rect 147 54 150 69
rect 3 39 6 49
rect 3 -8 6 34
rect 23 7 26 49
rect 42 24 45 49
rect 14 3 22 6
rect 23 -8 26 2
rect 42 -8 45 19
rect 55 -8 58 49
rect 74 24 77 49
rect 87 38 90 49
rect 74 -8 77 19
rect 87 -8 90 33
rect 102 17 105 49
rect 102 -8 105 12
rect 115 10 118 49
rect 137 12 140 49
rect 147 28 151 31
rect 115 -8 118 5
rect 137 -8 140 7
rect 14 -35 17 -16
rect 33 -35 36 -16
rect 65 -35 68 -16
rect 128 -35 131 -16
rect 147 -35 150 -16
rect -4 -37 157 -35
rect -4 -42 -2 -37
rect 3 -42 7 -37
rect 12 -42 17 -37
rect 22 -42 26 -37
rect 31 -42 35 -37
rect 40 -42 44 -37
rect 49 -42 53 -37
rect 58 -42 62 -37
rect 67 -42 72 -37
rect 77 -42 81 -37
rect 86 -42 91 -37
rect 96 -42 101 -37
rect 106 -42 111 -37
rect 116 -42 120 -37
rect 125 -42 130 -37
rect 135 -42 139 -37
rect 144 -42 148 -37
rect 153 -42 157 -37
rect -4 -46 157 -42
rect -4 -51 -2 -46
rect 3 -51 7 -46
rect 12 -51 17 -46
rect 22 -51 26 -46
rect 31 -51 35 -46
rect 40 -51 44 -46
rect 49 -51 53 -46
rect 58 -51 62 -46
rect 67 -51 72 -46
rect 77 -51 81 -46
rect 86 -51 91 -46
rect 96 -51 101 -46
rect 106 -51 111 -46
rect 116 -51 120 -46
rect 125 -51 130 -46
rect 135 -51 139 -46
rect 144 -51 148 -46
rect 153 -51 157 -46
rect -4 -53 157 -51
<< m2contact >>
rect 3 34 7 39
rect 48 27 52 32
rect 42 19 46 24
rect 29 12 33 17
rect 10 2 14 7
rect 22 2 26 7
rect 48 -2 52 3
rect 80 41 84 46
rect 86 33 90 38
rect 73 19 77 24
rect 61 5 65 10
rect 108 28 112 33
rect 101 12 105 17
rect 94 -6 98 -1
rect 122 19 126 24
rect 143 27 147 32
rect 115 5 119 10
rect 136 7 140 12
rect 108 -2 112 3
<< metal2 >>
rect 7 35 86 38
rect 46 19 73 22
rect 77 20 122 23
rect 33 13 101 16
rect -6 3 10 6
rect 65 6 115 9
<< m3contact >>
rect 80 41 84 46
rect 48 27 52 32
rect 108 28 112 33
rect 143 27 147 32
rect 136 7 140 12
rect 48 -2 52 3
rect 94 -6 98 -1
rect 108 -2 112 3
<< metal3 >>
rect 52 28 108 31
rect 112 28 143 31
rect 94 -1 97 28
<< m4contact >>
rect 80 41 84 46
rect 48 -2 52 3
rect 136 7 140 12
rect 108 -2 112 3
<< metal4 >>
rect 80 11 83 41
rect 80 8 136 11
rect 80 3 83 8
rect 52 0 83 3
rect 108 3 111 8
<< labels >>
rlabel metal1 70 -45 70 -45 1 vdd!
rlabel metal1 71 78 71 78 1 gnd!
rlabel metal1 151 28 151 31 1 clk
rlabel metal2 -6 3 -6 6 3 q
<< end >>
