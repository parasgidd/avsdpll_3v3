****************************
*PFD
***************************

.include osu018.lib


*______________________________________________
XX1 N001 N005 N002 VDD 0 nand101
XX2 N002 N008 N006 VDD 0 nand101
XX3 N006 N007 N008 VDD 0 nand101
XX4 N007 N010 N011 VDD 0 nand101
XX5 N011 N009 N010 VDD 0 nand101
XX6 N013 N012 N009 VDD 0 nand101
XX7 f_clk_in N005 VDD 0 inv101
XX8 f_VCO N013 VDD 0 inv101
XX9 N002 N003 VDD 0 inv101
XX10 N003 N004 VDD 0 inv101
XX11 N009 N014 VDD 0 inv101
XX12 N014 N015 VDD 0 inv101
XX13 N004 N006 N007 N001 VDD 0 nand301
XX14 N007 N010 N015 N012 VDD 0 nand301
XX15 N012 down VDD 0 inv101
XX16 N006 N002 N009 N010 VDD 0 N007 nand401
XX17 N001 up VDD 0 inv101



*______________________________________________
* _______SUBCIRCUITS_________________
*______________________________________________

.subckt nand101 in1 in2 out VDD GND
M1 out in1 N001 N001 nfet l=180n w=180n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 GND GND nfet l=180n w=360n
.ends nand101

.subckt inv101 in out VDD GND
M1 out in GND GND nfet l=180n w=180n
M2 VDD in out VDD pfet l=180n w=360n
.ends inv101

.subckt nand301 in1 in2 in3 out VDD GND
M1 out in1 N001 N001 nfet l=180n w=540n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 N002 N002 nfet l=180n w=540n
M5 N002 in3 GND GND nfet l=180n w=540n
M6 VDD in3 out VDD pfet l=180n w=360n
.ends nand301

.subckt nand401 in1 in2 in3 in4 VDD GND out
M1 out in1 N001 N001 nfet l=180n w=720n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 N002 N002 nfet l=180n w=720n
M5 N002 in3 N003 N003 nfet l=180n w=720n
M6 VDD in3 out VDD pfet l=180n w=360n
M7 N003 in4 GND GND nfet l=180n w=720n
M8 VDD in4 out VDD pfet l=180n w=360n
.ends nand401
*______________________________________________
* _______SUBCIRCUITS_ENDS________________
*______________________________________________


V1 f_clk_in 0 pulse 0 1.8 0 100p 100p 5n 10n
V2 f_VCO 0 pulse 0 1.8 2n 100p 100p 5n 9n
V3 VDD 0 1.8


.control
tran .1ns 50n
plot V(f_clk_in)+6 V(f_VCO)+4 V(up)+2 V(down)
.endc


.end
