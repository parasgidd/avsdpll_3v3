magic
tech scmos
timestamp 1599349060
<< nwell >>
rect 5 313 186 353
rect 52 293 186 313
rect 299 265 342 288
rect 251 235 342 265
rect 251 224 300 235
rect 52 117 124 140
rect 5 80 186 117
rect 349 8 374 154
rect 3 -133 491 -108
<< ntransistor >>
rect 16 411 18 414
rect 41 410 43 416
rect 51 410 53 416
rect 76 411 78 414
rect 100 411 102 414
rect 125 406 127 415
rect 136 406 138 415
rect 147 406 149 415
rect 173 411 175 414
rect 262 272 264 275
rect 278 272 280 275
rect 64 229 66 235
rect 74 229 76 235
rect 100 229 102 235
rect 110 229 112 235
rect 133 228 135 241
rect 139 228 141 241
rect 145 228 147 241
rect 151 228 153 241
rect 262 214 264 217
rect 278 214 280 217
rect 291 211 294 213
rect 318 212 321 214
rect 64 198 66 204
rect 74 198 76 204
rect 100 198 102 204
rect 110 198 112 204
rect 299 186 301 202
rect 311 199 313 202
rect 318 141 321 143
rect 318 125 321 127
rect 318 120 321 122
rect 318 104 321 106
rect 318 99 321 101
rect 16 19 18 22
rect 41 17 43 23
rect 51 17 53 23
rect 76 19 78 22
rect 100 19 102 22
rect 125 18 127 27
rect 136 18 138 27
rect 147 18 149 27
rect 318 83 321 85
rect 318 78 321 80
rect 318 62 321 64
rect 318 57 321 59
rect 318 41 321 43
rect 318 36 321 38
rect 173 19 175 22
rect 318 19 321 21
rect 17 -56 19 -53
rect 36 -56 38 -53
rect 56 -56 58 -53
rect 68 -56 70 -53
rect 86 -56 88 -53
rect 102 -56 104 -53
rect 116 -56 118 -53
rect 129 -56 131 -53
rect 150 -56 152 -53
rect 180 -56 182 -53
rect 199 -56 201 -53
rect 219 -56 221 -53
rect 231 -56 233 -53
rect 249 -56 251 -53
rect 265 -56 267 -53
rect 279 -56 281 -53
rect 292 -56 294 -53
rect 313 -56 315 -53
rect 343 -56 345 -53
rect 362 -56 364 -53
rect 382 -56 384 -53
rect 394 -56 396 -53
rect 412 -56 414 -53
rect 428 -56 430 -53
rect 442 -56 444 -53
rect 455 -56 457 -53
rect 476 -56 478 -53
<< ptransistor >>
rect 16 336 18 347
rect 41 336 43 347
rect 51 336 53 347
rect 76 336 78 347
rect 100 336 102 347
rect 125 336 127 347
rect 136 336 138 347
rect 147 336 149 347
rect 173 336 175 347
rect 64 299 66 310
rect 74 299 76 310
rect 100 299 102 310
rect 110 299 112 310
rect 133 299 135 310
rect 144 299 146 310
rect 155 299 157 310
rect 166 299 168 310
rect 262 251 264 259
rect 278 251 280 259
rect 294 251 296 259
rect 313 242 315 281
rect 329 261 336 263
rect 323 242 325 250
rect 262 230 264 238
rect 278 230 280 238
rect 355 141 361 143
rect 64 123 66 134
rect 74 123 76 134
rect 100 123 102 134
rect 110 123 112 134
rect 355 125 361 127
rect 355 120 361 122
rect 355 104 361 106
rect 355 99 361 101
rect 16 86 18 97
rect 41 86 43 97
rect 51 86 53 97
rect 76 86 78 97
rect 100 86 102 97
rect 125 86 127 97
rect 136 86 138 97
rect 147 86 149 97
rect 173 86 175 97
rect 355 83 361 85
rect 355 78 361 80
rect 355 62 361 64
rect 355 57 361 59
rect 355 41 361 43
rect 355 36 361 38
rect 355 19 361 21
rect 17 -122 19 -114
rect 36 -122 38 -114
rect 56 -122 58 -114
rect 68 -122 70 -114
rect 86 -122 88 -114
rect 102 -122 104 -114
rect 116 -122 118 -114
rect 129 -122 131 -114
rect 150 -122 152 -114
rect 180 -122 182 -114
rect 199 -122 201 -114
rect 219 -122 221 -114
rect 231 -122 233 -114
rect 249 -122 251 -114
rect 265 -122 267 -114
rect 279 -122 281 -114
rect 292 -122 294 -114
rect 313 -122 315 -114
rect 343 -122 345 -114
rect 362 -122 364 -114
rect 382 -122 384 -114
rect 394 -122 396 -114
rect 412 -122 414 -114
rect 428 -122 430 -114
rect 442 -122 444 -114
rect 455 -122 457 -114
rect 476 -122 478 -114
<< ndiffusion >>
rect 15 411 16 414
rect 18 411 19 414
rect 39 410 41 416
rect 43 410 51 416
rect 53 410 55 416
rect 75 411 76 414
rect 78 411 79 414
rect 99 411 100 414
rect 102 411 103 414
rect 123 406 125 415
rect 127 406 136 415
rect 138 406 147 415
rect 149 406 151 415
rect 172 411 173 414
rect 175 411 176 414
rect 261 272 262 275
rect 264 272 265 275
rect 277 272 278 275
rect 280 272 281 275
rect 62 229 64 235
rect 66 229 74 235
rect 76 229 78 235
rect 98 229 100 235
rect 102 229 110 235
rect 112 229 114 235
rect 131 228 133 241
rect 135 228 139 241
rect 141 228 145 241
rect 147 228 151 241
rect 153 228 159 241
rect 261 214 262 217
rect 264 214 265 217
rect 277 214 278 217
rect 280 214 281 217
rect 291 213 294 214
rect 318 214 321 219
rect 62 198 64 204
rect 66 198 74 204
rect 76 198 78 204
rect 98 198 100 204
rect 102 198 110 204
rect 112 198 114 204
rect 291 210 294 211
rect 318 210 321 212
rect 295 186 299 202
rect 301 186 305 202
rect 310 199 311 202
rect 313 199 314 202
rect 318 143 321 144
rect 318 140 321 141
rect 318 127 321 128
rect 318 122 321 125
rect 318 119 321 120
rect 318 106 321 107
rect 318 101 321 104
rect 318 98 321 99
rect 15 19 16 22
rect 18 19 19 22
rect 39 17 41 23
rect 43 17 51 23
rect 53 17 55 23
rect 75 19 76 22
rect 78 19 79 22
rect 99 19 100 22
rect 102 19 103 22
rect 123 18 125 27
rect 127 18 136 27
rect 138 18 147 27
rect 149 18 151 27
rect 318 85 321 86
rect 318 80 321 83
rect 318 77 321 78
rect 318 64 321 65
rect 318 59 321 62
rect 318 56 321 57
rect 318 43 321 44
rect 318 38 321 41
rect 318 35 321 36
rect 172 19 173 22
rect 175 19 176 22
rect 318 21 321 23
rect 318 18 321 19
rect 14 -56 17 -53
rect 19 -56 20 -53
rect 34 -56 36 -53
rect 38 -56 39 -53
rect 53 -56 56 -53
rect 58 -56 61 -53
rect 66 -56 68 -53
rect 70 -56 71 -53
rect 85 -56 86 -53
rect 88 -56 93 -53
rect 98 -56 102 -53
rect 104 -56 108 -53
rect 113 -56 116 -53
rect 118 -56 121 -53
rect 126 -56 129 -53
rect 131 -56 134 -53
rect 148 -56 150 -53
rect 152 -56 153 -53
rect 177 -56 180 -53
rect 182 -56 183 -53
rect 197 -56 199 -53
rect 201 -56 202 -53
rect 216 -56 219 -53
rect 221 -56 224 -53
rect 229 -56 231 -53
rect 233 -56 234 -53
rect 248 -56 249 -53
rect 251 -56 256 -53
rect 261 -56 265 -53
rect 267 -56 271 -53
rect 276 -56 279 -53
rect 281 -56 284 -53
rect 289 -56 292 -53
rect 294 -56 297 -53
rect 311 -56 313 -53
rect 315 -56 316 -53
rect 340 -56 343 -53
rect 345 -56 346 -53
rect 360 -56 362 -53
rect 364 -56 365 -53
rect 379 -56 382 -53
rect 384 -56 387 -53
rect 392 -56 394 -53
rect 396 -56 397 -53
rect 411 -56 412 -53
rect 414 -56 419 -53
rect 424 -56 428 -53
rect 430 -56 434 -53
rect 439 -56 442 -53
rect 444 -56 447 -53
rect 452 -56 455 -53
rect 457 -56 460 -53
rect 474 -56 476 -53
rect 478 -56 479 -53
<< pdiffusion >>
rect 15 336 16 347
rect 18 336 19 347
rect 39 336 41 347
rect 43 336 45 347
rect 49 336 51 347
rect 53 336 55 347
rect 75 336 76 347
rect 78 336 79 347
rect 99 336 100 347
rect 102 336 103 347
rect 123 336 125 347
rect 127 336 130 347
rect 134 336 136 347
rect 138 336 141 347
rect 145 336 147 347
rect 149 336 152 347
rect 172 336 173 347
rect 175 336 176 347
rect 62 299 64 310
rect 66 299 68 310
rect 72 299 74 310
rect 76 299 78 310
rect 98 299 100 310
rect 102 299 104 310
rect 108 299 110 310
rect 112 299 114 310
rect 131 299 133 310
rect 135 299 138 310
rect 142 299 144 310
rect 146 299 149 310
rect 153 299 155 310
rect 157 299 160 310
rect 164 299 166 310
rect 168 299 171 310
rect 261 251 262 259
rect 264 251 265 259
rect 277 251 278 259
rect 280 251 281 259
rect 293 251 294 259
rect 296 251 298 259
rect 310 242 313 281
rect 315 242 317 281
rect 329 263 336 266
rect 329 259 336 261
rect 321 242 323 250
rect 325 242 326 250
rect 261 230 262 238
rect 264 230 265 238
rect 277 230 278 238
rect 280 230 281 238
rect 355 143 361 144
rect 355 140 361 141
rect 62 123 64 134
rect 66 123 68 134
rect 72 123 74 134
rect 76 123 78 134
rect 98 123 100 134
rect 102 123 104 134
rect 108 123 110 134
rect 112 123 114 134
rect 355 127 361 128
rect 355 122 361 125
rect 355 119 361 120
rect 355 106 361 107
rect 355 101 361 104
rect 355 98 361 99
rect 15 86 16 97
rect 18 86 19 97
rect 39 86 41 97
rect 43 86 45 97
rect 49 86 51 97
rect 53 86 55 97
rect 75 86 76 97
rect 78 86 79 97
rect 99 86 100 97
rect 102 86 103 97
rect 123 86 125 97
rect 127 86 130 97
rect 134 86 136 97
rect 138 86 141 97
rect 145 86 147 97
rect 149 86 152 97
rect 172 86 173 97
rect 175 86 176 97
rect 355 85 361 86
rect 355 80 361 83
rect 355 77 361 78
rect 355 64 361 65
rect 355 59 361 62
rect 355 56 361 57
rect 355 43 361 44
rect 355 38 361 41
rect 355 35 361 36
rect 355 21 361 22
rect 355 18 361 19
rect 14 -122 17 -114
rect 19 -122 20 -114
rect 34 -122 36 -114
rect 38 -122 39 -114
rect 53 -122 56 -114
rect 58 -122 61 -114
rect 66 -122 68 -114
rect 70 -122 71 -114
rect 85 -122 86 -114
rect 88 -122 93 -114
rect 98 -122 102 -114
rect 104 -122 108 -114
rect 113 -122 116 -114
rect 118 -122 121 -114
rect 126 -122 129 -114
rect 131 -122 134 -114
rect 148 -122 150 -114
rect 152 -122 153 -114
rect 177 -122 180 -114
rect 182 -122 183 -114
rect 197 -122 199 -114
rect 201 -122 202 -114
rect 216 -122 219 -114
rect 221 -122 224 -114
rect 229 -122 231 -114
rect 233 -122 234 -114
rect 248 -122 249 -114
rect 251 -122 256 -114
rect 261 -122 265 -114
rect 267 -122 271 -114
rect 276 -122 279 -114
rect 281 -122 284 -114
rect 289 -122 292 -114
rect 294 -122 297 -114
rect 311 -122 313 -114
rect 315 -122 316 -114
rect 340 -122 343 -114
rect 345 -122 346 -114
rect 360 -122 362 -114
rect 364 -122 365 -114
rect 379 -122 382 -114
rect 384 -122 387 -114
rect 392 -122 394 -114
rect 396 -122 397 -114
rect 411 -122 412 -114
rect 414 -122 419 -114
rect 424 -122 428 -114
rect 430 -122 434 -114
rect 439 -122 442 -114
rect 444 -122 447 -114
rect 452 -122 455 -114
rect 457 -122 460 -114
rect 474 -122 476 -114
rect 478 -122 479 -114
<< ndcontact >>
rect 11 410 15 415
rect 19 410 23 415
rect 35 410 39 416
rect 55 410 59 416
rect 71 410 75 415
rect 79 410 83 415
rect 95 410 99 415
rect 103 410 107 415
rect 119 406 123 415
rect 151 406 155 415
rect 168 410 172 415
rect 176 410 180 415
rect 257 271 261 276
rect 265 271 269 276
rect 273 271 277 276
rect 281 271 285 276
rect 58 229 62 235
rect 78 229 82 235
rect 94 229 98 235
rect 114 229 118 235
rect 127 228 131 241
rect 159 228 163 241
rect 257 213 261 218
rect 265 213 269 218
rect 273 213 277 218
rect 317 219 322 223
rect 281 213 285 218
rect 290 214 295 218
rect 58 198 62 204
rect 78 198 82 204
rect 94 198 98 204
rect 114 198 118 204
rect 290 206 295 210
rect 317 206 322 210
rect 290 186 295 202
rect 305 186 310 202
rect 314 197 318 202
rect 317 144 322 148
rect 317 136 322 140
rect 317 128 322 132
rect 317 115 322 119
rect 317 107 322 111
rect 317 94 322 98
rect 317 86 322 90
rect 11 18 15 23
rect 19 18 23 23
rect 35 17 39 23
rect 55 17 59 23
rect 71 18 75 23
rect 79 18 83 23
rect 95 18 99 23
rect 103 18 107 23
rect 119 18 123 27
rect 151 18 155 27
rect 168 18 172 23
rect 317 73 322 77
rect 317 65 322 69
rect 317 52 322 56
rect 317 44 322 48
rect 317 31 322 35
rect 317 23 322 27
rect 176 18 180 23
rect 317 14 322 18
rect 9 -57 14 -52
rect 20 -57 25 -52
rect 29 -57 34 -52
rect 39 -57 44 -52
rect 48 -57 53 -52
rect 61 -57 66 -52
rect 71 -57 76 -52
rect 80 -57 85 -52
rect 93 -57 98 -52
rect 108 -57 113 -52
rect 121 -57 126 -52
rect 134 -57 139 -52
rect 143 -57 148 -52
rect 153 -57 158 -52
rect 172 -57 177 -52
rect 183 -57 188 -52
rect 192 -57 197 -52
rect 202 -57 207 -52
rect 211 -57 216 -52
rect 224 -57 229 -52
rect 234 -57 239 -52
rect 243 -57 248 -52
rect 256 -57 261 -52
rect 271 -57 276 -52
rect 284 -57 289 -52
rect 297 -57 302 -52
rect 306 -57 311 -52
rect 316 -57 321 -52
rect 335 -57 340 -52
rect 346 -57 351 -52
rect 355 -57 360 -52
rect 365 -57 370 -52
rect 374 -57 379 -52
rect 387 -57 392 -52
rect 397 -57 402 -52
rect 406 -57 411 -52
rect 419 -57 424 -52
rect 434 -57 439 -52
rect 447 -57 452 -52
rect 460 -57 465 -52
rect 469 -57 474 -52
rect 479 -57 484 -52
<< pdcontact >>
rect 11 336 15 347
rect 19 336 23 347
rect 35 336 39 347
rect 45 336 49 347
rect 55 336 59 347
rect 71 336 75 347
rect 79 336 83 347
rect 95 336 99 347
rect 103 336 107 347
rect 119 336 123 347
rect 130 336 134 347
rect 141 336 145 347
rect 152 336 156 347
rect 168 336 172 347
rect 176 336 180 347
rect 58 299 62 310
rect 68 299 72 310
rect 78 299 82 310
rect 94 299 98 310
rect 104 299 108 310
rect 114 299 118 310
rect 127 299 131 310
rect 138 299 142 310
rect 149 299 153 310
rect 160 299 164 310
rect 171 299 175 310
rect 257 251 261 259
rect 265 251 269 259
rect 273 251 277 259
rect 281 251 285 259
rect 289 251 293 259
rect 298 251 302 259
rect 306 242 310 281
rect 317 241 321 281
rect 329 266 336 270
rect 329 255 336 259
rect 326 242 330 250
rect 257 230 261 238
rect 265 230 269 238
rect 273 230 277 238
rect 281 230 285 238
rect 355 144 361 148
rect 355 136 361 140
rect 58 123 62 134
rect 68 123 72 134
rect 78 123 82 134
rect 94 123 98 134
rect 104 123 108 134
rect 114 123 118 134
rect 355 128 361 132
rect 355 115 361 119
rect 355 107 361 111
rect 11 86 15 97
rect 19 86 23 97
rect 35 86 39 97
rect 45 86 49 97
rect 55 86 59 97
rect 71 86 75 97
rect 79 86 83 97
rect 95 86 99 97
rect 103 86 107 97
rect 119 86 123 97
rect 130 86 134 97
rect 141 86 145 97
rect 152 86 156 97
rect 168 86 172 97
rect 176 86 180 97
rect 355 94 361 98
rect 355 86 361 90
rect 355 73 361 77
rect 355 65 361 69
rect 355 52 361 56
rect 355 44 361 48
rect 355 31 361 35
rect 355 22 361 26
rect 355 14 361 18
rect 9 -122 14 -114
rect 20 -122 25 -114
rect 29 -122 34 -114
rect 39 -122 44 -114
rect 48 -122 53 -114
rect 61 -122 66 -114
rect 71 -122 76 -114
rect 80 -122 85 -114
rect 93 -122 98 -114
rect 108 -122 113 -114
rect 121 -122 126 -114
rect 134 -122 139 -114
rect 143 -122 148 -114
rect 153 -122 158 -114
rect 172 -122 177 -114
rect 183 -122 188 -114
rect 192 -122 197 -114
rect 202 -122 207 -114
rect 211 -122 216 -114
rect 224 -122 229 -114
rect 234 -122 239 -114
rect 243 -122 248 -114
rect 256 -122 261 -114
rect 271 -122 276 -114
rect 284 -122 289 -114
rect 297 -122 302 -114
rect 306 -122 311 -114
rect 316 -122 321 -114
rect 335 -122 340 -114
rect 346 -122 351 -114
rect 355 -122 360 -114
rect 365 -122 370 -114
rect 374 -122 379 -114
rect 387 -122 392 -114
rect 397 -122 402 -114
rect 406 -122 411 -114
rect 419 -122 424 -114
rect 434 -122 439 -114
rect 447 -122 452 -114
rect 460 -122 465 -114
rect 469 -122 474 -114
rect 479 -122 484 -114
<< psubstratepcontact >>
rect 14 427 18 431
rect 22 427 26 431
rect 30 427 34 431
rect 38 427 42 431
rect 46 427 50 431
rect 54 427 58 431
rect 62 427 66 431
rect 70 427 74 431
rect 78 427 82 431
rect 86 427 90 431
rect 94 427 98 431
rect 102 427 106 431
rect 110 427 114 431
rect 118 427 122 431
rect 126 427 130 431
rect 134 427 138 431
rect 142 427 146 431
rect 150 427 154 431
rect 158 427 162 431
rect 166 427 170 431
rect 174 427 178 431
rect 182 427 186 431
rect 190 427 194 431
rect 198 427 202 431
rect 198 419 202 423
rect 198 411 202 415
rect 198 403 202 407
rect 198 395 202 399
rect 198 387 202 391
rect 198 379 202 383
rect 198 371 202 375
rect 198 363 202 367
rect 198 355 202 359
rect 198 342 202 346
rect 198 334 202 338
rect 198 325 202 329
rect 198 317 202 321
rect 198 309 202 313
rect 198 300 202 304
rect 198 292 202 296
rect 198 284 202 288
rect 198 276 202 280
rect 198 268 202 272
rect 198 260 202 264
rect 198 252 202 256
rect 198 244 202 248
rect 198 236 202 240
rect 198 228 202 232
rect 198 219 202 223
rect 58 214 62 218
rect 66 214 70 218
rect 74 214 78 218
rect 129 214 133 218
rect 137 214 141 218
rect 145 214 149 218
rect 154 214 158 218
rect 173 214 177 218
rect 181 214 185 218
rect 190 214 194 218
rect 198 211 202 215
rect 198 203 202 207
rect 198 195 202 199
rect 198 187 202 191
rect 198 179 202 183
rect 198 171 202 175
rect 198 163 202 167
rect 198 155 202 159
rect 198 147 202 151
rect 308 150 313 154
rect 198 138 202 142
rect 308 140 313 144
rect 198 130 202 134
rect 308 132 313 136
rect 198 122 202 126
rect 308 123 313 127
rect 198 114 202 118
rect 308 115 313 119
rect 198 106 202 110
rect 308 107 313 111
rect 198 98 202 102
rect 308 99 313 103
rect 198 90 202 94
rect 308 90 313 94
rect 198 82 202 86
rect 308 81 313 85
rect 198 74 202 78
rect 198 66 202 70
rect 308 66 313 70
rect 198 57 202 61
rect 308 58 313 62
rect 198 49 202 53
rect 308 50 313 54
rect 198 41 202 45
rect 308 40 313 44
rect 198 33 202 37
rect 308 32 313 36
rect 198 25 202 29
rect 308 24 313 28
rect 198 17 202 21
rect 308 16 313 20
rect 198 9 202 13
rect 308 8 313 12
rect 14 3 18 7
rect 22 3 26 7
rect 30 3 34 7
rect 38 3 42 7
rect 46 3 50 7
rect 54 3 58 7
rect 62 3 66 7
rect 70 3 74 7
rect 78 3 82 7
rect 86 3 90 7
rect 94 3 98 7
rect 102 3 106 7
rect 110 3 114 7
rect 118 3 122 7
rect 126 3 130 7
rect 134 3 138 7
rect 142 3 146 7
rect 150 3 154 7
rect 158 3 162 7
rect 166 3 170 7
rect 174 3 178 7
rect 182 3 186 7
rect 190 3 194 7
rect 198 1 202 5
rect 5 -26 10 -21
rect 14 -26 19 -21
rect 23 -26 28 -21
rect 32 -26 37 -21
rect 42 -26 47 -21
rect 51 -26 56 -21
rect 61 -26 66 -21
rect 70 -26 75 -21
rect 81 -26 86 -21
rect 91 -26 96 -21
rect 100 -26 105 -21
rect 109 -26 114 -21
rect 118 -26 123 -21
rect 127 -26 132 -21
rect 136 -26 141 -21
rect 145 -26 150 -21
rect 154 -26 159 -21
rect 168 -26 173 -21
rect 177 -26 182 -21
rect 186 -26 191 -21
rect 195 -26 200 -21
rect 205 -26 210 -21
rect 214 -26 219 -21
rect 224 -26 229 -21
rect 233 -26 238 -21
rect 244 -26 249 -21
rect 254 -26 259 -21
rect 263 -26 268 -21
rect 272 -26 277 -21
rect 281 -26 286 -21
rect 290 -26 295 -21
rect 299 -26 304 -21
rect 308 -26 313 -21
rect 317 -26 322 -21
rect 331 -26 336 -21
rect 340 -26 345 -21
rect 349 -26 354 -21
rect 358 -26 363 -21
rect 368 -26 373 -21
rect 377 -26 382 -21
rect 387 -26 392 -21
rect 396 -26 401 -21
rect 407 -26 412 -21
rect 417 -26 422 -21
rect 426 -26 431 -21
rect 435 -26 440 -21
rect 444 -26 449 -21
rect 453 -26 458 -21
rect 462 -26 467 -21
rect 471 -26 476 -21
rect 480 -26 485 -21
rect 5 -35 10 -30
rect 14 -35 19 -30
rect 23 -35 28 -30
rect 32 -35 37 -30
rect 42 -35 47 -30
rect 51 -35 56 -30
rect 61 -35 66 -30
rect 70 -35 75 -30
rect 81 -35 86 -30
rect 91 -35 96 -30
rect 100 -35 105 -30
rect 109 -35 114 -30
rect 118 -35 123 -30
rect 127 -35 132 -30
rect 136 -35 141 -30
rect 145 -35 150 -30
rect 154 -35 159 -30
rect 168 -35 173 -30
rect 177 -35 182 -30
rect 186 -35 191 -30
rect 195 -35 200 -30
rect 205 -35 210 -30
rect 214 -35 219 -30
rect 224 -35 229 -30
rect 233 -35 238 -30
rect 244 -35 249 -30
rect 254 -35 259 -30
rect 263 -35 268 -30
rect 272 -35 277 -30
rect 281 -35 286 -30
rect 290 -35 295 -30
rect 299 -35 304 -30
rect 308 -35 313 -30
rect 317 -35 322 -30
rect 331 -35 336 -30
rect 340 -35 345 -30
rect 349 -35 354 -30
rect 358 -35 363 -30
rect 368 -35 373 -30
rect 377 -35 382 -30
rect 387 -35 392 -30
rect 396 -35 401 -30
rect 407 -35 412 -30
rect 417 -35 422 -30
rect 426 -35 431 -30
rect 435 -35 440 -30
rect 444 -35 449 -30
rect 453 -35 458 -30
rect 462 -35 467 -30
rect 471 -35 476 -30
rect 480 -35 485 -30
<< nsubstratencontact >>
rect 8 325 12 329
rect 16 325 20 329
rect 26 325 30 329
rect 34 325 38 329
rect 51 325 55 329
rect 59 325 63 329
rect 119 325 123 329
rect 127 325 131 329
rect 137 325 141 329
rect 145 325 149 329
rect 8 317 12 321
rect 16 317 20 321
rect 26 317 30 321
rect 34 317 38 321
rect 51 317 55 321
rect 59 317 63 321
rect 119 317 123 321
rect 127 317 131 321
rect 137 317 141 321
rect 145 317 149 321
rect 366 147 371 151
rect 366 139 371 143
rect 366 131 371 135
rect 366 123 371 127
rect 366 115 371 119
rect 8 107 12 111
rect 16 107 20 111
rect 24 107 28 111
rect 32 107 36 111
rect 40 107 44 111
rect 49 107 53 111
rect 57 107 61 111
rect 117 108 121 112
rect 125 108 129 112
rect 133 108 137 112
rect 141 108 145 112
rect 149 108 153 112
rect 167 108 171 112
rect 366 107 371 111
rect 366 99 371 103
rect 366 91 371 95
rect 366 83 371 87
rect 366 75 371 79
rect 366 67 371 71
rect 366 59 371 63
rect 366 51 371 55
rect 366 43 371 47
rect 366 35 371 39
rect 366 27 371 31
rect 366 19 371 23
rect 366 11 371 15
rect 5 -148 10 -143
rect 14 -148 19 -143
rect 24 -148 29 -143
rect 33 -148 38 -143
rect 42 -148 47 -143
rect 51 -148 56 -143
rect 60 -148 65 -143
rect 69 -148 74 -143
rect 79 -148 84 -143
rect 88 -148 93 -143
rect 98 -148 103 -143
rect 108 -148 113 -143
rect 118 -148 123 -143
rect 127 -148 132 -143
rect 137 -148 142 -143
rect 146 -148 151 -143
rect 155 -148 160 -143
rect 168 -148 173 -143
rect 177 -148 182 -143
rect 187 -148 192 -143
rect 196 -148 201 -143
rect 205 -148 210 -143
rect 214 -148 219 -143
rect 223 -148 228 -143
rect 232 -148 237 -143
rect 242 -148 247 -143
rect 251 -148 256 -143
rect 261 -148 266 -143
rect 271 -148 276 -143
rect 281 -148 286 -143
rect 290 -148 295 -143
rect 300 -148 305 -143
rect 309 -148 314 -143
rect 318 -148 323 -143
rect 331 -148 336 -143
rect 340 -148 345 -143
rect 350 -148 355 -143
rect 359 -148 364 -143
rect 368 -148 373 -143
rect 377 -148 382 -143
rect 386 -148 391 -143
rect 395 -148 400 -143
rect 405 -148 410 -143
rect 414 -148 419 -143
rect 424 -148 429 -143
rect 434 -148 439 -143
rect 444 -148 449 -143
rect 453 -148 458 -143
rect 463 -148 468 -143
rect 472 -148 477 -143
rect 481 -148 486 -143
rect 5 -157 10 -152
rect 14 -157 19 -152
rect 24 -157 29 -152
rect 33 -157 38 -152
rect 42 -157 47 -152
rect 51 -157 56 -152
rect 60 -157 65 -152
rect 69 -157 74 -152
rect 79 -157 84 -152
rect 88 -157 93 -152
rect 98 -157 103 -152
rect 108 -157 113 -152
rect 118 -157 123 -152
rect 127 -157 132 -152
rect 137 -157 142 -152
rect 146 -157 151 -152
rect 155 -157 160 -152
rect 168 -157 173 -152
rect 177 -157 182 -152
rect 187 -157 192 -152
rect 196 -157 201 -152
rect 205 -157 210 -152
rect 214 -157 219 -152
rect 223 -157 228 -152
rect 232 -157 237 -152
rect 242 -157 247 -152
rect 251 -157 256 -152
rect 261 -157 266 -152
rect 271 -157 276 -152
rect 281 -157 286 -152
rect 290 -157 295 -152
rect 300 -157 305 -152
rect 309 -157 314 -152
rect 318 -157 323 -152
rect 331 -157 336 -152
rect 340 -157 345 -152
rect 350 -157 355 -152
rect 359 -157 364 -152
rect 368 -157 373 -152
rect 377 -157 382 -152
rect 386 -157 391 -152
rect 395 -157 400 -152
rect 405 -157 410 -152
rect 414 -157 419 -152
rect 424 -157 429 -152
rect 434 -157 439 -152
rect 444 -157 449 -152
rect 453 -157 458 -152
rect 463 -157 468 -152
rect 472 -157 477 -152
rect 481 -157 486 -152
<< polysilicon >>
rect 41 416 43 418
rect 51 416 53 418
rect 16 414 18 416
rect 16 347 18 411
rect 76 414 78 416
rect 41 347 43 410
rect 51 397 53 410
rect 52 392 53 397
rect 51 347 53 392
rect 76 347 78 411
rect 100 414 102 416
rect 125 415 127 417
rect 136 415 138 417
rect 147 415 149 417
rect 100 347 102 411
rect 173 414 175 416
rect 125 371 127 406
rect 125 347 127 366
rect 136 347 138 406
rect 147 377 149 406
rect 147 347 149 372
rect 173 347 175 411
rect 16 334 18 336
rect 41 334 43 336
rect 51 334 53 336
rect 76 334 78 336
rect 100 334 102 336
rect 125 334 127 336
rect 136 334 138 336
rect 147 334 149 336
rect 173 334 175 336
rect 64 310 66 312
rect 74 310 76 312
rect 100 310 102 312
rect 110 310 112 312
rect 133 310 135 312
rect 144 310 146 312
rect 155 310 157 312
rect 166 310 168 312
rect 64 235 66 299
rect 74 291 76 299
rect 74 235 76 286
rect 100 273 102 299
rect 100 235 102 268
rect 110 235 112 299
rect 133 273 135 299
rect 133 241 135 268
rect 144 265 146 299
rect 155 276 157 299
rect 143 263 146 265
rect 139 241 141 260
rect 155 252 157 271
rect 145 250 157 252
rect 145 241 147 250
rect 166 249 168 299
rect 279 279 280 283
rect 313 281 315 286
rect 262 275 264 277
rect 262 268 264 272
rect 278 275 280 279
rect 278 270 280 272
rect 263 264 264 268
rect 262 259 264 264
rect 278 259 280 261
rect 294 259 296 263
rect 262 249 264 251
rect 151 244 166 246
rect 278 246 280 251
rect 294 249 296 251
rect 151 241 153 244
rect 64 227 66 229
rect 74 227 76 229
rect 100 227 102 229
rect 110 227 112 229
rect 262 238 264 240
rect 278 238 280 241
rect 313 240 315 242
rect 324 263 326 273
rect 323 261 329 263
rect 336 261 338 263
rect 323 250 325 261
rect 323 240 325 242
rect 133 226 135 228
rect 139 226 141 228
rect 145 226 147 228
rect 151 226 153 228
rect 262 217 264 230
rect 278 228 280 230
rect 279 221 280 225
rect 262 210 264 214
rect 278 217 280 221
rect 278 212 280 214
rect 286 211 291 213
rect 294 211 296 213
rect 314 212 318 214
rect 321 212 323 214
rect 64 204 66 206
rect 74 204 76 206
rect 100 204 102 206
rect 110 204 112 206
rect 286 209 288 211
rect 285 205 288 209
rect 299 202 301 205
rect 311 202 313 212
rect 64 189 66 198
rect 64 134 66 184
rect 74 147 76 198
rect 100 164 102 198
rect 74 134 76 142
rect 100 134 102 160
rect 110 134 112 198
rect 311 197 313 199
rect 299 183 301 186
rect 316 141 318 143
rect 321 142 325 143
rect 321 141 330 142
rect 352 141 355 143
rect 361 141 363 143
rect 64 121 66 123
rect 74 121 76 123
rect 100 121 102 123
rect 110 121 112 123
rect 316 125 318 127
rect 321 126 325 127
rect 321 125 330 126
rect 352 125 355 127
rect 361 125 363 127
rect 316 120 318 122
rect 321 121 334 122
rect 339 121 355 122
rect 321 120 355 121
rect 361 120 363 122
rect 316 104 318 106
rect 321 105 325 106
rect 321 104 330 105
rect 352 104 355 106
rect 361 104 363 106
rect 16 97 18 99
rect 41 97 43 99
rect 51 97 53 99
rect 76 97 78 99
rect 100 97 102 99
rect 125 97 127 99
rect 136 97 138 99
rect 147 97 149 99
rect 173 97 175 99
rect 316 99 318 101
rect 321 100 333 101
rect 338 100 355 101
rect 321 99 355 100
rect 361 99 363 101
rect 16 22 18 86
rect 41 23 43 86
rect 51 41 53 86
rect 52 36 53 41
rect 51 23 53 36
rect 16 17 18 19
rect 76 22 78 86
rect 76 17 78 19
rect 100 22 102 86
rect 125 67 127 86
rect 125 27 127 62
rect 136 27 138 86
rect 147 61 149 86
rect 147 27 149 56
rect 100 17 102 19
rect 173 22 175 86
rect 316 83 318 85
rect 321 84 325 85
rect 321 83 330 84
rect 352 83 355 85
rect 361 83 363 85
rect 316 78 318 80
rect 321 79 333 80
rect 338 79 355 80
rect 321 78 355 79
rect 361 78 363 80
rect 316 62 318 64
rect 321 63 325 64
rect 321 62 330 63
rect 352 62 355 64
rect 361 62 363 64
rect 316 57 318 59
rect 321 58 333 59
rect 338 58 355 59
rect 321 57 355 58
rect 361 57 363 59
rect 316 41 318 43
rect 321 42 325 43
rect 321 41 330 42
rect 352 41 355 43
rect 361 41 363 43
rect 316 36 318 38
rect 321 37 333 38
rect 338 37 355 38
rect 321 36 355 37
rect 361 36 363 38
rect 41 15 43 17
rect 51 15 53 17
rect 125 16 127 18
rect 136 16 138 18
rect 147 16 149 18
rect 173 17 175 19
rect 316 19 318 21
rect 321 20 334 21
rect 339 20 355 21
rect 321 19 355 20
rect 361 19 363 21
rect 17 -53 19 -51
rect 17 -99 19 -56
rect 36 -53 38 -51
rect 36 -89 38 -56
rect 56 -53 58 -51
rect 56 -74 58 -56
rect 68 -53 70 -51
rect 17 -114 19 -104
rect 36 -114 38 -94
rect 68 -96 70 -56
rect 86 -53 88 -51
rect 86 -58 88 -56
rect 102 -53 104 -51
rect 102 -58 104 -56
rect 116 -53 118 -51
rect 86 -60 104 -58
rect 116 -73 118 -56
rect 129 -53 131 -51
rect 129 -82 131 -56
rect 150 -53 152 -51
rect 150 -74 152 -56
rect 180 -53 182 -51
rect 56 -114 58 -108
rect 68 -114 70 -101
rect 86 -112 101 -110
rect 86 -114 88 -112
rect 102 -114 104 -112
rect 116 -114 118 -108
rect 129 -114 131 -87
rect 150 -114 152 -79
rect 180 -99 182 -56
rect 199 -53 201 -51
rect 199 -89 201 -56
rect 219 -53 221 -51
rect 219 -74 221 -56
rect 231 -53 233 -51
rect 180 -114 182 -104
rect 199 -114 201 -94
rect 231 -96 233 -56
rect 249 -53 251 -51
rect 249 -58 251 -56
rect 265 -53 267 -51
rect 265 -58 267 -56
rect 279 -53 281 -51
rect 249 -60 267 -58
rect 279 -73 281 -56
rect 292 -53 294 -51
rect 292 -82 294 -56
rect 313 -53 315 -51
rect 313 -74 315 -56
rect 343 -53 345 -51
rect 219 -114 221 -108
rect 231 -114 233 -101
rect 249 -112 264 -110
rect 249 -114 251 -112
rect 265 -114 267 -112
rect 279 -114 281 -108
rect 292 -114 294 -87
rect 313 -114 315 -79
rect 343 -99 345 -56
rect 362 -53 364 -51
rect 362 -89 364 -56
rect 382 -53 384 -51
rect 382 -74 384 -56
rect 394 -53 396 -51
rect 343 -114 345 -104
rect 362 -114 364 -94
rect 394 -96 396 -56
rect 412 -53 414 -51
rect 412 -58 414 -56
rect 428 -53 430 -51
rect 428 -58 430 -56
rect 442 -53 444 -51
rect 412 -60 430 -58
rect 442 -73 444 -56
rect 455 -53 457 -51
rect 455 -82 457 -56
rect 476 -53 478 -51
rect 476 -74 478 -56
rect 382 -114 384 -108
rect 394 -114 396 -101
rect 412 -112 427 -110
rect 412 -114 414 -112
rect 428 -114 430 -112
rect 442 -114 444 -108
rect 455 -114 457 -87
rect 476 -114 478 -79
rect 17 -124 19 -122
rect 36 -124 38 -122
rect 56 -124 58 -122
rect 68 -124 70 -122
rect 86 -124 88 -122
rect 102 -124 104 -122
rect 116 -124 118 -122
rect 129 -124 131 -122
rect 150 -124 152 -122
rect 180 -124 182 -122
rect 199 -124 201 -122
rect 219 -124 221 -122
rect 231 -124 233 -122
rect 249 -124 251 -122
rect 265 -124 267 -122
rect 279 -124 281 -122
rect 292 -124 294 -122
rect 313 -124 315 -122
rect 343 -124 345 -122
rect 362 -124 364 -122
rect 382 -124 384 -122
rect 394 -124 396 -122
rect 412 -124 414 -122
rect 428 -124 430 -122
rect 442 -124 444 -122
rect 455 -124 457 -122
rect 476 -124 478 -122
<< polycontact >>
rect 11 378 16 383
rect 36 402 41 407
rect 48 392 52 397
rect 71 366 76 371
rect 53 356 58 361
rect 95 377 100 382
rect 132 377 136 382
rect 124 366 128 371
rect 168 399 173 404
rect 146 372 150 377
rect 60 271 64 276
rect 74 286 78 291
rect 98 268 102 273
rect 112 288 116 293
rect 131 268 135 273
rect 153 271 157 276
rect 139 260 143 265
rect 311 286 316 290
rect 274 279 279 283
rect 258 264 263 268
rect 293 263 297 268
rect 166 244 170 249
rect 277 241 281 246
rect 324 273 328 278
rect 274 221 279 225
rect 310 212 314 217
rect 261 206 266 210
rect 281 205 285 209
rect 63 184 67 189
rect 60 157 64 162
rect 97 160 102 164
rect 74 142 78 147
rect 112 176 117 180
rect 297 179 302 183
rect 325 142 330 146
rect 347 139 352 143
rect 325 126 330 130
rect 347 125 352 129
rect 334 121 339 125
rect 325 105 330 109
rect 347 104 352 108
rect 333 100 338 104
rect 11 50 16 55
rect 36 26 41 31
rect 53 72 58 77
rect 71 62 76 67
rect 48 36 52 41
rect 95 51 100 56
rect 124 62 128 67
rect 132 51 136 56
rect 146 56 150 61
rect 168 29 173 34
rect 325 84 330 88
rect 347 83 352 87
rect 333 79 338 83
rect 325 63 330 67
rect 347 62 352 66
rect 333 58 338 62
rect 325 42 330 46
rect 347 41 352 45
rect 333 37 338 41
rect 334 20 339 24
rect 55 -79 59 -74
rect 36 -94 40 -89
rect 17 -104 21 -99
rect 87 -65 91 -60
rect 115 -78 119 -73
rect 150 -79 154 -74
rect 129 -87 133 -82
rect 68 -101 72 -96
rect 55 -108 59 -103
rect 101 -112 105 -107
rect 115 -108 119 -103
rect 218 -79 222 -74
rect 199 -94 203 -89
rect 180 -104 184 -99
rect 250 -65 254 -60
rect 278 -78 282 -73
rect 313 -79 317 -74
rect 292 -87 296 -82
rect 231 -101 235 -96
rect 218 -108 222 -103
rect 264 -112 268 -107
rect 278 -108 282 -103
rect 381 -79 385 -74
rect 362 -94 366 -89
rect 343 -104 347 -99
rect 413 -65 417 -60
rect 441 -78 445 -73
rect 476 -79 480 -74
rect 455 -87 459 -82
rect 394 -101 398 -96
rect 381 -108 385 -103
rect 427 -112 431 -107
rect 441 -108 445 -103
<< metal1 >>
rect 11 431 205 434
rect 11 427 14 431
rect 18 427 22 431
rect 26 427 30 431
rect 34 427 38 431
rect 42 427 46 431
rect 50 427 54 431
rect 58 427 62 431
rect 66 427 70 431
rect 74 427 78 431
rect 82 427 86 431
rect 90 427 94 431
rect 98 427 102 431
rect 106 427 110 431
rect 114 427 118 431
rect 122 427 126 431
rect 130 427 134 431
rect 138 427 142 431
rect 146 427 150 431
rect 154 427 158 431
rect 162 427 166 431
rect 170 427 174 431
rect 178 427 182 431
rect 186 427 190 431
rect 194 427 198 431
rect 202 427 205 431
rect 11 424 205 427
rect 11 415 14 424
rect 35 416 38 424
rect 71 415 74 424
rect 95 415 98 424
rect 119 415 122 424
rect 168 415 171 424
rect 195 423 205 424
rect 195 419 198 423
rect 202 419 205 423
rect 195 415 205 419
rect 20 406 23 410
rect 20 403 36 406
rect 3 379 11 382
rect 20 347 23 403
rect 56 370 59 410
rect 80 381 83 410
rect 80 378 95 381
rect 45 367 71 370
rect 45 347 48 367
rect 80 347 83 378
rect 104 370 107 410
rect 152 403 155 406
rect 140 400 168 403
rect 140 396 143 400
rect 121 393 143 396
rect 104 367 124 370
rect 104 347 107 367
rect 140 360 143 393
rect 177 395 180 410
rect 195 411 198 415
rect 202 411 205 415
rect 195 407 205 411
rect 195 403 198 407
rect 202 403 205 407
rect 195 399 205 403
rect 177 392 186 395
rect 134 357 156 360
rect 130 347 133 356
rect 153 347 156 357
rect 177 347 180 392
rect 195 395 198 399
rect 202 395 205 399
rect 195 391 205 395
rect 11 330 14 336
rect 35 330 38 336
rect 56 330 59 336
rect 195 387 198 391
rect 202 387 205 391
rect 195 383 205 387
rect 195 379 198 383
rect 202 379 205 383
rect 195 375 205 379
rect 195 371 198 375
rect 202 371 205 375
rect 195 367 205 371
rect 195 363 198 367
rect 202 363 205 367
rect 195 359 205 363
rect 195 355 198 359
rect 202 355 205 359
rect 195 346 205 355
rect 195 342 198 346
rect 202 342 205 346
rect 195 338 205 342
rect 71 330 74 336
rect 95 330 98 336
rect 119 330 122 336
rect 141 330 144 336
rect 168 330 171 336
rect 195 334 198 338
rect 202 334 205 338
rect 5 329 175 330
rect 5 325 8 329
rect 12 325 16 329
rect 20 325 26 329
rect 30 325 34 329
rect 38 325 51 329
rect 55 325 59 329
rect 63 325 119 329
rect 123 325 127 329
rect 131 325 137 329
rect 141 325 145 329
rect 149 327 175 329
rect 149 325 168 327
rect 5 321 168 325
rect 5 317 8 321
rect 12 317 16 321
rect 20 317 26 321
rect 30 317 34 321
rect 38 317 51 321
rect 55 317 59 321
rect 63 317 119 321
rect 123 317 127 321
rect 131 317 137 321
rect 141 317 145 321
rect 149 317 168 321
rect 5 316 168 317
rect 5 117 23 316
rect 58 310 61 316
rect 79 310 82 316
rect 94 310 97 316
rect 115 310 118 316
rect 127 310 130 316
rect 149 310 152 316
rect 172 310 175 316
rect 195 329 205 334
rect 195 325 198 329
rect 202 325 205 329
rect 195 321 205 325
rect 195 317 198 321
rect 202 317 205 321
rect 195 313 205 317
rect 195 309 198 313
rect 202 309 205 313
rect 195 304 205 309
rect 195 300 198 304
rect 202 300 205 304
rect 68 279 71 299
rect 104 290 107 299
rect 78 287 107 290
rect 138 292 141 299
rect 116 289 141 292
rect 104 284 107 287
rect 138 287 141 289
rect 160 287 163 299
rect 138 284 163 287
rect 104 281 118 284
rect 68 276 82 279
rect 79 272 82 276
rect 79 269 98 272
rect 79 235 82 269
rect 115 235 118 281
rect 160 241 163 284
rect 195 296 205 300
rect 195 292 198 296
rect 202 292 205 296
rect 195 288 205 292
rect 195 284 198 288
rect 202 284 205 288
rect 195 283 205 284
rect 282 286 311 289
rect 195 280 248 283
rect 195 276 198 280
rect 202 279 248 280
rect 202 276 205 279
rect 282 276 285 286
rect 195 272 205 276
rect 195 268 198 272
rect 202 268 205 272
rect 269 273 273 276
rect 195 264 205 268
rect 195 260 198 264
rect 202 260 205 264
rect 195 256 205 260
rect 266 259 269 271
rect 282 259 285 271
rect 195 252 198 256
rect 202 252 205 256
rect 195 248 205 252
rect 269 256 273 259
rect 195 244 198 248
rect 202 244 205 248
rect 58 223 61 229
rect 94 223 97 229
rect 195 240 205 244
rect 195 236 198 240
rect 202 236 205 240
rect 195 232 205 236
rect 195 228 198 232
rect 202 228 205 232
rect 269 230 273 233
rect 127 223 130 228
rect 195 223 205 228
rect 58 219 198 223
rect 202 219 205 223
rect 58 218 205 219
rect 266 218 269 230
rect 282 218 285 230
rect 327 228 330 242
rect 327 225 337 228
rect 313 220 317 223
rect 62 214 66 218
rect 70 214 74 218
rect 78 214 129 218
rect 133 214 137 218
rect 141 214 145 218
rect 149 214 154 218
rect 158 214 173 218
rect 177 214 181 218
rect 185 214 190 218
rect 194 217 205 218
rect 194 215 247 217
rect 194 214 198 215
rect 58 211 198 214
rect 202 212 247 215
rect 269 213 273 216
rect 295 215 302 218
rect 202 211 205 212
rect 58 209 205 211
rect 58 204 61 209
rect 94 204 97 209
rect 195 207 205 209
rect 195 203 198 207
rect 202 203 205 207
rect 282 209 285 213
rect 266 206 276 209
rect 79 164 82 198
rect 115 194 118 198
rect 195 199 205 203
rect 195 195 198 199
rect 202 195 205 199
rect 105 191 118 194
rect 79 161 97 164
rect 79 157 82 161
rect 68 154 82 157
rect 68 134 71 154
rect 105 152 108 191
rect 160 179 163 195
rect 195 191 205 195
rect 195 187 198 191
rect 202 187 205 191
rect 195 183 205 187
rect 117 176 163 179
rect 195 179 198 183
rect 202 179 205 183
rect 273 182 276 206
rect 299 209 302 215
rect 310 217 313 220
rect 295 206 308 209
rect 305 202 308 206
rect 327 202 330 225
rect 318 199 330 202
rect 104 149 108 152
rect 160 151 163 176
rect 104 146 107 149
rect 78 143 107 146
rect 104 134 107 143
rect 58 117 61 123
rect 79 117 82 123
rect 94 117 97 123
rect 115 117 118 123
rect 5 112 171 117
rect 5 111 117 112
rect 5 107 8 111
rect 12 107 16 111
rect 20 107 24 111
rect 28 107 32 111
rect 36 107 40 111
rect 44 107 49 111
rect 53 107 57 111
rect 61 108 117 111
rect 121 108 125 112
rect 129 108 133 112
rect 137 108 141 112
rect 145 108 149 112
rect 153 108 167 112
rect 61 107 171 108
rect 5 103 171 107
rect 11 97 14 103
rect 35 97 38 103
rect 56 97 59 103
rect 71 97 74 103
rect 95 97 98 103
rect 119 97 122 103
rect 141 97 144 103
rect 168 97 171 103
rect 177 97 180 176
rect -10 51 11 54
rect -10 -98 -5 51
rect 20 30 23 86
rect 45 66 48 86
rect 45 63 71 66
rect 20 27 36 30
rect 20 23 23 27
rect 56 23 59 63
rect 80 55 83 86
rect 104 66 107 86
rect 130 77 133 86
rect 153 76 156 86
rect 134 73 156 76
rect 104 63 124 66
rect 80 52 95 55
rect 80 23 83 52
rect 104 23 107 63
rect 140 40 143 73
rect 121 37 143 40
rect 140 33 143 37
rect 177 41 180 86
rect 195 175 205 179
rect 277 179 297 182
rect 195 171 198 175
rect 202 171 205 175
rect 195 167 205 171
rect 195 163 198 167
rect 202 163 205 167
rect 195 159 205 163
rect 195 155 198 159
rect 202 155 205 159
rect 195 151 205 155
rect 195 147 198 151
rect 202 147 205 151
rect 195 142 205 147
rect 195 138 198 142
rect 202 138 205 142
rect 195 134 205 138
rect 195 130 198 134
rect 202 130 205 134
rect 195 126 205 130
rect 195 122 198 126
rect 202 122 205 126
rect 195 118 205 122
rect 195 114 198 118
rect 202 114 205 118
rect 195 110 205 114
rect 195 106 198 110
rect 202 106 205 110
rect 195 102 205 106
rect 195 98 198 102
rect 202 98 205 102
rect 195 94 205 98
rect 195 90 198 94
rect 202 90 205 94
rect 195 86 205 90
rect 195 82 198 86
rect 202 82 205 86
rect 195 78 205 82
rect 195 74 198 78
rect 202 74 205 78
rect 195 70 205 74
rect 195 66 198 70
rect 202 66 205 70
rect 195 61 205 66
rect 195 57 198 61
rect 202 57 205 61
rect 195 53 205 57
rect 195 49 198 53
rect 202 49 205 53
rect 195 45 205 49
rect 195 41 198 45
rect 202 41 205 45
rect 177 38 185 41
rect 140 30 168 33
rect 152 27 155 30
rect 11 10 14 18
rect 177 23 180 38
rect 195 37 205 41
rect 195 33 198 37
rect 202 33 205 37
rect 195 29 205 33
rect 195 25 198 29
rect 202 25 205 29
rect 195 21 205 25
rect 35 10 38 17
rect 71 10 74 18
rect 95 10 98 18
rect 119 10 122 18
rect 168 10 171 18
rect 195 17 198 21
rect 202 17 205 21
rect 195 13 205 17
rect 195 10 198 13
rect 11 9 198 10
rect 202 9 205 13
rect 11 7 205 9
rect 308 148 313 150
rect 308 145 317 148
rect 308 144 313 145
rect 325 146 330 199
rect 366 151 374 154
rect 361 147 366 148
rect 371 147 374 151
rect 361 145 374 147
rect 366 143 374 145
rect 308 136 313 140
rect 322 136 355 139
rect 371 139 374 143
rect 366 135 374 139
rect 308 129 317 132
rect 308 127 313 129
rect 361 131 366 132
rect 371 131 374 135
rect 361 129 374 131
rect 366 127 374 129
rect 308 119 313 123
rect 371 123 374 127
rect 366 119 374 123
rect 322 115 355 118
rect 371 115 374 119
rect 308 111 313 115
rect 313 108 317 111
rect 308 103 313 107
rect 333 104 336 115
rect 366 111 374 115
rect 361 108 366 111
rect 371 107 374 111
rect 366 103 374 107
rect 308 94 313 99
rect 371 99 374 103
rect 322 94 355 97
rect 366 95 374 99
rect 308 87 317 90
rect 308 85 313 87
rect 308 70 313 81
rect 333 83 336 94
rect 371 91 374 95
rect 366 90 374 91
rect 361 87 374 90
rect 371 83 374 87
rect 366 79 374 83
rect 322 73 355 76
rect 371 75 374 79
rect 313 66 317 69
rect 308 62 313 66
rect 333 62 336 73
rect 366 71 374 75
rect 361 67 366 69
rect 371 67 374 71
rect 361 66 374 67
rect 366 63 374 66
rect 371 59 374 63
rect 308 54 313 58
rect 322 52 355 55
rect 366 55 374 59
rect 308 48 313 50
rect 308 45 317 48
rect 308 44 313 45
rect 308 36 313 40
rect 333 41 336 52
rect 371 51 374 55
rect 366 48 374 51
rect 361 47 374 48
rect 361 45 366 47
rect 371 43 374 47
rect 366 39 374 43
rect 371 35 374 39
rect 308 28 313 32
rect 322 31 334 34
rect 339 31 355 34
rect 366 31 374 35
rect 313 24 317 27
rect 308 20 313 24
rect 334 24 339 30
rect 371 27 374 31
rect 366 26 374 27
rect 361 23 374 26
rect 371 19 374 23
rect 308 12 313 16
rect 322 14 355 17
rect 366 15 374 19
rect 11 3 14 7
rect 18 3 22 7
rect 26 3 30 7
rect 34 3 38 7
rect 42 3 46 7
rect 50 3 54 7
rect 58 3 62 7
rect 66 3 70 7
rect 74 3 78 7
rect 82 3 86 7
rect 90 3 94 7
rect 98 3 102 7
rect 106 3 110 7
rect 114 3 118 7
rect 122 3 126 7
rect 130 3 134 7
rect 138 3 142 7
rect 146 3 150 7
rect 154 3 158 7
rect 162 3 166 7
rect 170 3 174 7
rect 178 3 182 7
rect 186 3 190 7
rect 194 5 205 7
rect 194 3 198 5
rect 11 1 198 3
rect 202 1 205 5
rect 11 0 205 1
rect 334 2 339 14
rect 371 11 374 15
rect 366 8 374 11
rect 334 -3 504 2
rect 3 -21 490 -17
rect 3 -26 5 -21
rect 10 -26 14 -21
rect 19 -26 23 -21
rect 28 -26 32 -21
rect 37 -26 42 -21
rect 47 -26 51 -21
rect 56 -26 61 -21
rect 66 -26 70 -21
rect 75 -26 81 -21
rect 86 -26 91 -21
rect 96 -26 100 -21
rect 105 -26 109 -21
rect 114 -26 118 -21
rect 123 -26 127 -21
rect 132 -26 136 -21
rect 141 -26 145 -21
rect 150 -26 154 -21
rect 159 -26 168 -21
rect 173 -26 177 -21
rect 182 -26 186 -21
rect 191 -26 195 -21
rect 200 -26 205 -21
rect 210 -26 214 -21
rect 219 -26 224 -21
rect 229 -26 233 -21
rect 238 -26 244 -21
rect 249 -26 254 -21
rect 259 -26 263 -21
rect 268 -26 272 -21
rect 277 -26 281 -21
rect 286 -26 290 -21
rect 295 -26 299 -21
rect 304 -26 308 -21
rect 313 -26 317 -21
rect 322 -26 331 -21
rect 336 -26 340 -21
rect 345 -26 349 -21
rect 354 -26 358 -21
rect 363 -26 368 -21
rect 373 -26 377 -21
rect 382 -26 387 -21
rect 392 -26 396 -21
rect 401 -26 407 -21
rect 412 -26 417 -21
rect 422 -26 426 -21
rect 431 -26 435 -21
rect 440 -26 444 -21
rect 449 -26 453 -21
rect 458 -26 462 -21
rect 467 -26 471 -21
rect 476 -26 480 -21
rect 485 -26 490 -21
rect 3 -30 490 -26
rect 3 -35 5 -30
rect 10 -35 14 -30
rect 19 -35 23 -30
rect 28 -35 32 -30
rect 37 -35 42 -30
rect 47 -35 51 -30
rect 56 -35 61 -30
rect 66 -35 70 -30
rect 75 -35 81 -30
rect 86 -35 91 -30
rect 96 -35 100 -30
rect 105 -35 109 -30
rect 114 -35 118 -30
rect 123 -35 127 -30
rect 132 -35 136 -30
rect 141 -35 145 -30
rect 150 -35 154 -30
rect 159 -35 168 -30
rect 173 -35 177 -30
rect 182 -35 186 -30
rect 191 -35 195 -30
rect 200 -35 205 -30
rect 210 -35 214 -30
rect 219 -35 224 -30
rect 229 -35 233 -30
rect 238 -35 244 -30
rect 249 -35 254 -30
rect 259 -35 263 -30
rect 268 -35 272 -30
rect 277 -35 281 -30
rect 286 -35 290 -30
rect 295 -35 299 -30
rect 304 -35 308 -30
rect 313 -35 317 -30
rect 322 -35 331 -30
rect 336 -35 340 -30
rect 345 -35 349 -30
rect 354 -35 358 -30
rect 363 -35 368 -30
rect 373 -35 377 -30
rect 382 -35 387 -30
rect 392 -35 396 -30
rect 401 -35 407 -30
rect 412 -35 417 -30
rect 422 -35 426 -30
rect 431 -35 435 -30
rect 440 -35 444 -30
rect 449 -35 453 -30
rect 458 -35 462 -30
rect 467 -35 471 -30
rect 476 -35 480 -30
rect 485 -35 490 -30
rect 3 -37 490 -35
rect 21 -52 24 -37
rect 40 -52 43 -37
rect 72 -52 75 -37
rect 135 -52 138 -37
rect 154 -52 157 -37
rect 184 -52 187 -37
rect 203 -52 206 -37
rect 235 -52 238 -37
rect 298 -52 301 -37
rect 317 -52 320 -37
rect 347 -52 350 -37
rect 366 -52 369 -37
rect 398 -52 401 -37
rect 461 -52 464 -37
rect 480 -52 483 -37
rect 10 -67 13 -57
rect 10 -114 13 -72
rect 30 -99 33 -57
rect 49 -82 52 -57
rect 21 -103 29 -100
rect 30 -114 33 -104
rect 49 -114 52 -87
rect 62 -114 65 -57
rect 81 -82 84 -57
rect 94 -68 97 -57
rect 81 -114 84 -87
rect 94 -114 97 -73
rect 109 -89 112 -57
rect 109 -114 112 -94
rect 122 -96 125 -57
rect 144 -94 147 -57
rect 173 -67 176 -57
rect 154 -78 161 -75
rect 122 -114 125 -101
rect 144 -114 147 -99
rect 173 -114 176 -72
rect 193 -99 196 -57
rect 212 -82 215 -57
rect 184 -103 192 -100
rect 193 -114 196 -104
rect 212 -114 215 -87
rect 225 -114 228 -57
rect 244 -82 247 -57
rect 257 -68 260 -57
rect 244 -114 247 -87
rect 257 -114 260 -73
rect 272 -89 275 -57
rect 272 -114 275 -94
rect 285 -96 288 -57
rect 307 -94 310 -57
rect 336 -67 339 -57
rect 317 -78 324 -75
rect 285 -114 288 -101
rect 307 -114 310 -99
rect 336 -114 339 -72
rect 356 -99 359 -57
rect 375 -82 378 -57
rect 347 -103 355 -100
rect 356 -114 359 -104
rect 375 -114 378 -87
rect 388 -114 391 -57
rect 407 -82 410 -57
rect 420 -68 423 -57
rect 407 -114 410 -87
rect 420 -114 423 -73
rect 435 -89 438 -57
rect 435 -114 438 -94
rect 448 -96 451 -57
rect 470 -94 473 -57
rect 499 -75 504 -3
rect 480 -78 504 -75
rect 448 -114 451 -101
rect 470 -114 473 -99
rect 21 -141 24 -122
rect 40 -141 43 -122
rect 72 -141 75 -122
rect 135 -141 138 -122
rect 154 -141 157 -122
rect 184 -141 187 -122
rect 203 -141 206 -122
rect 235 -141 238 -122
rect 298 -141 301 -122
rect 317 -141 320 -122
rect 347 -141 350 -122
rect 366 -141 369 -122
rect 398 -141 401 -122
rect 461 -141 464 -122
rect 480 -141 483 -122
rect 3 -143 490 -141
rect 3 -148 5 -143
rect 10 -148 14 -143
rect 19 -148 24 -143
rect 29 -148 33 -143
rect 38 -148 42 -143
rect 47 -148 51 -143
rect 56 -148 60 -143
rect 65 -148 69 -143
rect 74 -148 79 -143
rect 84 -148 88 -143
rect 93 -148 98 -143
rect 103 -148 108 -143
rect 113 -148 118 -143
rect 123 -148 127 -143
rect 132 -148 137 -143
rect 142 -148 146 -143
rect 151 -148 155 -143
rect 160 -148 168 -143
rect 173 -148 177 -143
rect 182 -148 187 -143
rect 192 -148 196 -143
rect 201 -148 205 -143
rect 210 -148 214 -143
rect 219 -148 223 -143
rect 228 -148 232 -143
rect 237 -148 242 -143
rect 247 -148 251 -143
rect 256 -148 261 -143
rect 266 -148 271 -143
rect 276 -148 281 -143
rect 286 -148 290 -143
rect 295 -148 300 -143
rect 305 -148 309 -143
rect 314 -148 318 -143
rect 323 -148 331 -143
rect 336 -148 340 -143
rect 345 -148 350 -143
rect 355 -148 359 -143
rect 364 -148 368 -143
rect 373 -148 377 -143
rect 382 -148 386 -143
rect 391 -148 395 -143
rect 400 -148 405 -143
rect 410 -148 414 -143
rect 419 -148 424 -143
rect 429 -148 434 -143
rect 439 -148 444 -143
rect 449 -148 453 -143
rect 458 -148 463 -143
rect 468 -148 472 -143
rect 477 -148 481 -143
rect 486 -148 490 -143
rect 3 -152 490 -148
rect 3 -157 5 -152
rect 10 -157 14 -152
rect 19 -157 24 -152
rect 29 -157 33 -152
rect 38 -157 42 -152
rect 47 -157 51 -152
rect 56 -157 60 -152
rect 65 -157 69 -152
rect 74 -157 79 -152
rect 84 -157 88 -152
rect 93 -157 98 -152
rect 103 -157 108 -152
rect 113 -157 118 -152
rect 123 -157 127 -152
rect 132 -157 137 -152
rect 142 -157 146 -152
rect 151 -157 155 -152
rect 160 -157 168 -152
rect 173 -157 177 -152
rect 182 -157 187 -152
rect 192 -157 196 -152
rect 201 -157 205 -152
rect 210 -157 214 -152
rect 219 -157 223 -152
rect 228 -157 232 -152
rect 237 -157 242 -152
rect 247 -157 251 -152
rect 256 -157 261 -152
rect 266 -157 271 -152
rect 276 -157 281 -152
rect 286 -157 290 -152
rect 295 -157 300 -152
rect 305 -157 309 -152
rect 314 -157 318 -152
rect 323 -157 331 -152
rect 336 -157 340 -152
rect 345 -157 350 -152
rect 355 -157 359 -152
rect 364 -157 368 -152
rect 373 -157 377 -152
rect 382 -157 386 -152
rect 391 -157 395 -152
rect 400 -157 405 -152
rect 410 -157 414 -152
rect 419 -157 424 -152
rect 429 -157 434 -152
rect 439 -157 444 -152
rect 449 -157 453 -152
rect 458 -157 463 -152
rect 468 -157 472 -152
rect 477 -157 481 -152
rect 486 -157 490 -152
rect 3 -159 490 -157
<< m2contact >>
rect 48 392 52 397
rect 53 356 58 361
rect 117 392 121 397
rect 132 377 136 382
rect 129 356 134 361
rect 146 372 150 377
rect 186 391 190 396
rect 45 336 49 347
rect 168 316 175 327
rect 68 299 72 310
rect 160 299 164 310
rect 60 271 64 276
rect 98 268 102 273
rect 131 268 135 273
rect 153 271 157 276
rect 139 260 143 265
rect 248 279 253 283
rect 274 279 279 283
rect 257 271 261 276
rect 258 264 263 268
rect 293 263 297 268
rect 166 244 170 249
rect 257 251 261 259
rect 289 251 293 259
rect 298 251 302 259
rect 159 228 163 241
rect 277 241 281 246
rect 306 242 310 252
rect 324 273 328 278
rect 329 266 336 270
rect 317 255 321 260
rect 329 255 336 259
rect 274 221 279 225
rect 307 220 313 224
rect 247 212 253 217
rect 257 213 261 218
rect 78 198 82 204
rect 63 184 67 189
rect 159 195 164 200
rect 60 157 64 162
rect 176 176 181 182
rect 317 206 322 210
rect 290 186 295 202
rect 159 146 164 151
rect 68 123 72 134
rect 45 86 49 97
rect 53 72 58 77
rect 48 36 52 41
rect 129 72 134 77
rect 132 51 136 56
rect 117 36 121 41
rect 146 56 150 61
rect 272 177 277 182
rect 325 142 330 146
rect 347 139 352 143
rect 325 126 330 130
rect 347 125 352 129
rect 334 121 339 125
rect 325 105 330 109
rect 347 104 352 108
rect 325 84 330 88
rect 347 83 352 87
rect 325 63 330 67
rect 347 62 352 66
rect 325 42 330 46
rect 347 41 352 45
rect 334 30 339 34
rect -10 -103 -5 -98
rect 10 -72 14 -67
rect 55 -79 59 -74
rect 49 -87 53 -82
rect 36 -94 40 -89
rect 17 -104 21 -99
rect 29 -104 33 -99
rect 55 -108 59 -103
rect 87 -65 91 -60
rect 93 -73 97 -68
rect 80 -87 84 -82
rect 68 -101 72 -96
rect 115 -78 119 -73
rect 108 -94 112 -89
rect 101 -112 105 -107
rect 129 -87 133 -82
rect 173 -72 177 -67
rect 150 -79 154 -74
rect 161 -80 165 -75
rect 122 -101 126 -96
rect 143 -99 147 -94
rect 115 -108 119 -103
rect 218 -79 222 -74
rect 212 -87 216 -82
rect 199 -94 203 -89
rect 180 -104 184 -99
rect 192 -104 196 -99
rect 218 -108 222 -103
rect 250 -65 254 -60
rect 256 -73 260 -68
rect 243 -87 247 -82
rect 231 -101 235 -96
rect 278 -78 282 -73
rect 271 -94 275 -89
rect 264 -112 268 -107
rect 292 -87 296 -82
rect 336 -72 340 -67
rect 313 -79 317 -74
rect 324 -80 328 -75
rect 285 -101 289 -96
rect 306 -99 310 -94
rect 278 -108 282 -103
rect 381 -79 385 -74
rect 375 -87 379 -82
rect 362 -94 366 -89
rect 343 -104 347 -99
rect 355 -104 359 -99
rect 381 -108 385 -103
rect 413 -65 417 -60
rect 419 -73 423 -68
rect 406 -87 410 -82
rect 394 -101 398 -96
rect 441 -78 445 -73
rect 434 -94 438 -89
rect 427 -112 431 -107
rect 455 -87 459 -82
rect 476 -79 480 -74
rect 448 -101 452 -96
rect 469 -99 473 -94
rect 441 -108 445 -103
<< metal2 >>
rect 190 391 245 396
rect 58 357 129 360
rect 160 310 163 376
rect 102 269 131 272
rect 240 267 245 391
rect 253 280 274 283
rect 253 279 260 280
rect 279 280 328 283
rect 257 276 260 279
rect 324 278 328 280
rect 328 273 334 276
rect 331 270 334 273
rect 240 264 258 267
rect 263 264 293 267
rect 302 256 317 259
rect 289 246 292 251
rect 299 246 302 251
rect 289 243 302 246
rect 181 178 272 182
rect 325 130 330 142
rect 58 73 129 76
rect 160 57 163 117
rect 325 109 330 126
rect 347 129 352 139
rect 325 88 330 105
rect 325 67 330 84
rect 325 46 330 63
rect 347 108 352 125
rect 347 87 352 104
rect 347 66 352 83
rect 347 45 352 62
rect 14 -71 93 -68
rect 177 -71 256 -68
rect 340 -71 419 -68
rect 53 -87 80 -84
rect 84 -86 129 -83
rect 40 -93 108 -90
rect -5 -103 17 -100
rect 72 -100 122 -97
rect 162 -100 165 -80
rect 216 -87 243 -84
rect 247 -86 292 -83
rect 203 -93 271 -90
rect 162 -103 180 -100
rect 235 -100 285 -97
rect 325 -100 328 -80
rect 379 -87 406 -84
rect 410 -86 455 -83
rect 366 -93 434 -90
rect 325 -103 343 -100
rect 398 -100 448 -97
<< m3contact >>
rect 48 392 52 397
rect 117 392 121 397
rect 132 377 136 382
rect 146 372 150 377
rect 45 336 49 347
rect 168 316 175 327
rect 68 299 72 310
rect 160 299 164 310
rect 60 271 64 276
rect 153 271 157 276
rect 139 260 143 265
rect 257 251 261 259
rect 329 255 336 259
rect 166 244 170 249
rect 277 241 281 246
rect 306 242 310 252
rect 159 228 163 241
rect 274 221 279 225
rect 307 220 313 224
rect 247 212 253 217
rect 257 213 261 218
rect 317 206 322 210
rect 78 198 82 204
rect 159 195 164 200
rect 63 184 67 189
rect 290 186 295 202
rect 60 157 64 162
rect 159 146 164 151
rect 68 123 72 134
rect 45 86 49 97
rect 146 56 150 61
rect 334 121 339 125
rect 132 51 136 56
rect 48 36 52 41
rect 117 36 121 41
rect 334 30 339 34
rect 87 -65 91 -60
rect 250 -65 254 -60
rect 413 -65 417 -60
rect 55 -79 59 -74
rect 115 -78 119 -73
rect 150 -79 154 -74
rect 218 -79 222 -74
rect 278 -78 282 -73
rect 313 -79 317 -74
rect 381 -79 385 -74
rect 441 -78 445 -73
rect 476 -79 480 -74
rect 143 -99 147 -94
rect 55 -108 59 -103
rect 101 -112 105 -107
rect 115 -108 119 -103
rect 306 -99 310 -94
rect 218 -108 222 -103
rect 264 -112 268 -107
rect 278 -108 282 -103
rect 469 -99 473 -94
rect 381 -108 385 -103
rect 427 -112 431 -107
rect 441 -108 445 -103
<< metal3 >>
rect 52 393 117 396
rect 112 378 132 381
rect 45 275 48 336
rect 112 323 115 378
rect 150 373 163 376
rect 68 320 115 323
rect 68 310 71 320
rect 160 310 163 373
rect 168 327 233 328
rect 175 316 233 327
rect 45 272 60 275
rect 64 272 153 275
rect 121 262 139 265
rect 121 218 124 262
rect 223 249 233 316
rect 257 249 261 251
rect 223 246 306 249
rect 223 245 261 246
rect 79 215 124 218
rect 79 204 82 215
rect 160 200 163 228
rect 167 188 170 244
rect 257 230 261 245
rect 331 249 334 255
rect 310 246 334 249
rect 257 221 274 224
rect 307 224 310 242
rect 279 221 295 224
rect 257 218 260 221
rect 253 213 257 216
rect 292 209 295 221
rect 292 206 317 209
rect 292 202 295 206
rect 67 184 170 188
rect 45 158 60 161
rect 45 97 48 158
rect 68 113 71 123
rect 68 110 115 113
rect 112 55 115 110
rect 160 60 163 146
rect 150 57 163 60
rect 112 52 132 55
rect 52 37 117 40
rect 59 -78 115 -75
rect 119 -78 150 -75
rect 101 -107 104 -78
rect 222 -78 278 -75
rect 282 -78 313 -75
rect 264 -107 267 -78
rect 385 -78 441 -75
rect 445 -78 476 -75
rect 427 -107 430 -78
<< m4contact >>
rect 334 121 339 125
rect 334 30 339 34
rect 87 -65 91 -60
rect 250 -65 254 -60
rect 413 -65 417 -60
rect 55 -108 59 -103
rect 143 -99 147 -94
rect 115 -108 119 -103
rect 218 -108 222 -103
rect 306 -99 310 -94
rect 278 -108 282 -103
rect 381 -108 385 -103
rect 469 -99 473 -94
rect 441 -108 445 -103
<< metal4 >>
rect 334 34 339 121
rect 87 -95 90 -65
rect 87 -98 143 -95
rect 87 -103 90 -98
rect 59 -106 90 -103
rect 115 -103 118 -98
rect 250 -95 253 -65
rect 250 -98 306 -95
rect 250 -103 253 -98
rect 222 -106 253 -103
rect 278 -103 281 -98
rect 413 -95 416 -65
rect 413 -98 469 -95
rect 413 -103 416 -98
rect 385 -106 416 -103
rect 441 -103 444 -98
<< labels >>
rlabel metal1 3 379 3 382 3 fin
rlabel metal1 3 51 3 54 3 fvco_8
rlabel metal1 185 38 185 41 1 dn
rlabel metal1 200 216 200 216 7 gnd!
rlabel metal1 14 218 14 218 1 vdd!
rlabel metal1 185 392 185 395 1 up
rlabel metal1 337 225 337 228 7 cp
rlabel metal1 78 -28 78 -28 1 gnd!
rlabel metal1 241 -28 241 -28 1 gnd!
rlabel metal1 404 -28 404 -28 1 gnd!
rlabel metal1 403 -151 403 -151 1 vdd!
rlabel metal1 240 -151 240 -151 1 vdd!
rlabel metal1 77 -151 77 -151 1 vdd!
rlabel metal1 334 8 339 8 1 fout
rlabel metal1 372 81 372 81 7 vdd!
rlabel metal1 311 78 311 78 3 gnd!
<< end >>
