magic
tech scmos
timestamp 1598605816
<< nwell >>
rect -2 52 140 93
rect -2 -96 140 -55
<< ntransistor >>
rect 10 128 12 131
rect 28 128 30 131
rect 36 128 38 131
rect 52 128 54 131
rect 69 128 71 131
rect 86 128 88 131
rect 91 128 93 131
rect 96 128 98 131
rect 122 128 124 131
rect 48 5 50 8
rect 56 5 58 8
rect 75 5 77 8
rect 83 5 85 8
rect 103 5 105 8
rect 108 5 110 8
rect 113 5 115 8
rect 118 5 120 8
rect 48 -22 50 -19
rect 56 -22 58 -19
rect 75 -22 77 -19
rect 83 -22 85 -19
rect 10 -135 12 -132
rect 28 -135 30 -132
rect 36 -135 38 -132
rect 52 -135 54 -132
rect 69 -135 71 -132
rect 86 -135 88 -132
rect 91 -135 93 -132
rect 96 -135 98 -132
rect 122 -135 124 -132
<< ptransistor >>
rect 10 79 12 87
rect 28 79 30 87
rect 36 79 38 87
rect 52 79 54 87
rect 69 79 71 87
rect 86 79 88 87
rect 94 79 96 87
rect 102 79 104 87
rect 122 79 124 87
rect 48 58 50 66
rect 56 58 58 66
rect 75 58 77 66
rect 83 58 85 66
rect 103 58 105 66
rect 111 58 113 66
rect 119 58 121 66
rect 127 58 129 66
rect 48 -69 50 -61
rect 56 -69 58 -61
rect 75 -69 77 -61
rect 83 -69 85 -61
rect 10 -90 12 -82
rect 28 -90 30 -82
rect 36 -90 38 -82
rect 52 -90 54 -82
rect 69 -90 71 -82
rect 86 -90 88 -82
rect 94 -90 96 -82
rect 102 -90 104 -82
rect 122 -90 124 -82
<< ndiffusion >>
rect 9 128 10 131
rect 12 128 14 131
rect 27 128 28 131
rect 30 128 36 131
rect 38 128 39 131
rect 51 128 52 131
rect 54 128 56 131
rect 68 128 69 131
rect 71 128 73 131
rect 85 128 86 131
rect 88 128 91 131
rect 93 128 96 131
rect 98 128 100 131
rect 104 128 111 131
rect 121 128 122 131
rect 124 128 126 131
rect 47 5 48 8
rect 50 5 56 8
rect 58 5 59 8
rect 74 5 75 8
rect 77 5 83 8
rect 85 5 86 8
rect 102 5 103 8
rect 105 5 108 8
rect 110 5 113 8
rect 115 5 118 8
rect 120 5 121 8
rect 47 -22 48 -19
rect 50 -22 56 -19
rect 58 -22 59 -19
rect 74 -22 75 -19
rect 77 -22 83 -19
rect 85 -22 86 -19
rect 9 -135 10 -132
rect 12 -135 14 -132
rect 27 -135 28 -132
rect 30 -135 36 -132
rect 38 -135 39 -132
rect 51 -135 52 -132
rect 54 -135 56 -132
rect 68 -135 69 -132
rect 71 -135 73 -132
rect 85 -135 86 -132
rect 88 -135 91 -132
rect 93 -135 96 -132
rect 98 -135 100 -132
rect 104 -135 111 -132
rect 121 -135 122 -132
rect 124 -135 126 -132
<< pdiffusion >>
rect 9 79 10 87
rect 12 79 14 87
rect 27 79 28 87
rect 30 79 31 87
rect 35 79 36 87
rect 38 79 39 87
rect 51 79 52 87
rect 54 79 56 87
rect 68 79 69 87
rect 71 79 73 87
rect 85 79 86 87
rect 88 79 89 87
rect 93 79 94 87
rect 96 79 97 87
rect 101 79 102 87
rect 104 79 105 87
rect 109 79 110 87
rect 121 79 122 87
rect 124 79 126 87
rect 47 58 48 66
rect 50 58 51 66
rect 55 58 56 66
rect 58 58 59 66
rect 74 58 75 66
rect 77 58 78 66
rect 82 58 83 66
rect 85 58 86 66
rect 102 58 103 66
rect 105 58 106 66
rect 110 58 111 66
rect 113 58 114 66
rect 118 58 119 66
rect 121 58 122 66
rect 126 58 127 66
rect 129 58 130 66
rect 47 -69 48 -61
rect 50 -69 51 -61
rect 55 -69 56 -61
rect 58 -69 59 -61
rect 74 -69 75 -61
rect 77 -69 78 -61
rect 82 -69 83 -61
rect 85 -69 86 -61
rect 9 -90 10 -82
rect 12 -90 14 -82
rect 27 -90 28 -82
rect 30 -90 31 -82
rect 35 -90 36 -82
rect 38 -90 39 -82
rect 51 -90 52 -82
rect 54 -90 56 -82
rect 68 -90 69 -82
rect 71 -90 73 -82
rect 85 -90 86 -82
rect 88 -90 89 -82
rect 93 -90 94 -82
rect 96 -90 97 -82
rect 101 -90 102 -82
rect 104 -90 105 -82
rect 109 -90 110 -82
rect 121 -90 122 -82
rect 124 -90 126 -82
<< ndcontact >>
rect 5 127 9 132
rect 14 127 18 132
rect 23 127 27 132
rect 39 127 43 132
rect 47 127 51 132
rect 56 127 60 132
rect 64 127 68 132
rect 73 127 77 132
rect 81 127 85 132
rect 100 127 104 132
rect 117 127 121 132
rect 126 127 130 132
rect 43 4 47 9
rect 59 4 63 9
rect 70 4 74 9
rect 86 4 90 9
rect 98 4 102 9
rect 121 4 125 9
rect 43 -23 47 -18
rect 59 -23 63 -18
rect 70 -23 74 -18
rect 86 -23 90 -18
rect 5 -136 9 -131
rect 14 -136 18 -131
rect 23 -136 27 -131
rect 39 -136 43 -131
rect 47 -136 51 -131
rect 56 -136 60 -131
rect 64 -136 68 -131
rect 73 -136 77 -131
rect 81 -136 85 -131
rect 100 -136 104 -131
rect 117 -136 121 -131
rect 126 -136 130 -131
<< pdcontact >>
rect 5 79 9 87
rect 14 79 18 87
rect 23 79 27 87
rect 31 79 35 87
rect 39 79 43 87
rect 47 79 51 87
rect 56 79 60 87
rect 64 79 68 87
rect 73 79 77 87
rect 81 79 85 87
rect 89 79 93 87
rect 97 79 101 87
rect 105 79 109 87
rect 117 79 121 87
rect 126 79 130 87
rect 43 58 47 66
rect 51 58 55 66
rect 59 58 63 66
rect 70 58 74 66
rect 78 58 82 66
rect 86 58 90 66
rect 98 58 102 66
rect 106 58 110 66
rect 114 58 118 66
rect 122 58 126 66
rect 130 58 134 66
rect 43 -69 47 -61
rect 51 -69 55 -61
rect 59 -69 63 -61
rect 70 -69 74 -61
rect 78 -69 82 -61
rect 86 -69 90 -61
rect 5 -90 9 -82
rect 14 -90 18 -82
rect 23 -90 27 -82
rect 31 -90 35 -82
rect 39 -90 43 -82
rect 47 -90 51 -82
rect 56 -90 60 -82
rect 64 -90 68 -82
rect 73 -90 77 -82
rect 81 -90 85 -82
rect 89 -90 93 -82
rect 97 -90 101 -82
rect 105 -90 109 -82
rect 117 -90 121 -82
rect 126 -90 130 -82
<< psubstratepcontact >>
rect 0 139 5 144
rect 9 139 14 144
rect 18 139 23 144
rect 27 139 32 144
rect 36 139 41 144
rect 45 139 50 144
rect 54 139 59 144
rect 63 139 68 144
rect 72 139 77 144
rect 81 139 86 144
rect 90 139 95 144
rect 99 139 104 144
rect 108 139 113 144
rect 117 139 122 144
rect 126 139 131 144
rect 135 139 140 144
rect 149 137 154 142
rect 149 128 154 133
rect 149 118 154 123
rect 149 108 154 113
rect 149 96 154 101
rect 149 84 154 89
rect 149 75 154 80
rect 149 65 154 70
rect 149 54 154 59
rect 149 45 154 50
rect 149 36 154 41
rect 149 27 154 32
rect 149 18 154 23
rect 149 9 154 14
rect 149 0 154 5
rect 40 -10 45 -5
rect 49 -10 54 -5
rect 58 -10 63 -5
rect 67 -10 72 -5
rect 76 -10 81 -5
rect 85 -10 90 -5
rect 94 -10 99 -5
rect 103 -10 108 -5
rect 113 -10 118 -5
rect 140 -10 145 -5
rect 149 -11 154 -6
rect 148 -23 153 -18
rect 148 -35 153 -30
rect 148 -46 153 -41
rect 148 -57 153 -52
rect 148 -68 153 -63
rect 148 -78 153 -73
rect 148 -89 153 -84
rect 148 -99 153 -94
rect 148 -109 153 -104
rect 148 -119 153 -114
rect 148 -128 153 -123
rect 148 -137 153 -132
rect 0 -148 5 -143
rect 9 -148 14 -143
rect 18 -148 23 -143
rect 27 -148 32 -143
rect 36 -148 41 -143
rect 45 -148 50 -143
rect 54 -148 59 -143
rect 63 -148 68 -143
rect 72 -148 77 -143
rect 81 -148 86 -143
rect 90 -148 95 -143
rect 99 -148 104 -143
rect 108 -148 113 -143
rect 117 -148 122 -143
rect 126 -148 131 -143
rect 135 -148 140 -143
rect 148 -148 153 -143
<< nsubstratencontact >>
rect 38 70 43 75
rect 47 70 52 75
rect 56 70 61 75
rect 65 70 70 75
rect 74 70 79 75
rect 83 70 88 75
rect 92 70 97 75
rect 101 70 106 75
rect 110 70 115 75
rect 119 70 124 75
rect 128 70 133 75
rect 1 64 6 69
rect 10 64 15 69
rect 19 64 24 69
rect 1 55 6 60
rect 10 55 15 60
rect 19 55 24 60
rect 1 44 6 49
rect 1 34 6 39
rect 1 25 6 30
rect 1 16 6 21
rect 1 7 6 12
rect 1 -2 6 3
rect 1 -11 6 -6
rect 1 -20 6 -15
rect 1 -30 6 -25
rect 1 -40 6 -35
rect 1 -53 6 -48
rect 1 -63 6 -58
rect 10 -63 15 -58
rect 19 -63 24 -58
rect 119 -69 124 -64
rect 128 -69 133 -64
rect 1 -74 6 -69
rect 10 -74 15 -69
rect 19 -74 24 -69
rect 28 -78 33 -73
rect 38 -78 43 -73
rect 47 -78 52 -73
rect 56 -78 61 -73
rect 65 -78 70 -73
rect 74 -78 79 -73
rect 83 -78 88 -73
rect 92 -78 97 -73
rect 101 -78 106 -73
rect 110 -78 115 -73
rect 119 -78 124 -73
rect 128 -78 133 -73
<< polysilicon >>
rect 10 131 12 133
rect 10 100 12 128
rect 28 131 30 133
rect 36 131 38 133
rect 28 111 30 128
rect 36 107 38 128
rect 52 131 54 133
rect 52 118 54 128
rect 69 131 71 133
rect 69 123 71 128
rect 86 131 88 133
rect 91 131 93 133
rect 96 131 98 133
rect 10 87 12 96
rect 28 87 30 107
rect 36 87 38 102
rect 52 87 54 113
rect 69 87 71 119
rect 86 106 88 128
rect 91 113 93 128
rect 96 118 98 128
rect 122 131 124 133
rect 96 116 104 118
rect 86 87 88 101
rect 94 87 96 108
rect 102 106 104 116
rect 102 103 107 106
rect 102 87 104 103
rect 122 98 124 128
rect 122 87 124 94
rect 10 77 12 79
rect 28 77 30 79
rect 36 77 38 79
rect 52 77 54 79
rect 69 77 71 79
rect 86 77 88 79
rect 94 77 96 79
rect 102 77 104 79
rect 122 77 124 79
rect 48 66 50 68
rect 56 66 58 68
rect 75 66 77 68
rect 83 66 85 68
rect 103 66 105 68
rect 111 66 113 68
rect 119 66 121 68
rect 127 66 129 68
rect 48 48 50 58
rect 48 8 50 44
rect 56 38 58 58
rect 56 8 58 33
rect 75 31 77 58
rect 83 27 85 58
rect 48 3 50 5
rect 56 3 58 5
rect 75 8 77 26
rect 84 22 85 27
rect 83 8 85 22
rect 75 3 77 5
rect 83 3 85 5
rect 103 8 105 58
rect 111 44 113 58
rect 108 8 110 40
rect 119 34 121 58
rect 118 32 121 34
rect 113 8 115 30
rect 127 17 129 58
rect 123 15 129 17
rect 118 8 120 14
rect 103 3 105 5
rect 108 3 110 5
rect 113 3 115 5
rect 118 3 120 5
rect 48 -19 50 -17
rect 56 -19 58 -17
rect 48 -26 50 -22
rect 48 -47 50 -31
rect 48 -61 50 -51
rect 56 -43 58 -22
rect 75 -19 77 -17
rect 83 -19 85 -17
rect 75 -36 77 -22
rect 83 -31 85 -22
rect 84 -36 85 -31
rect 56 -61 58 -48
rect 75 -61 77 -41
rect 83 -61 85 -36
rect 48 -71 50 -69
rect 56 -71 58 -69
rect 75 -71 77 -69
rect 83 -71 85 -69
rect 10 -82 12 -80
rect 28 -82 30 -80
rect 36 -82 38 -80
rect 52 -82 54 -80
rect 69 -82 71 -80
rect 86 -82 88 -80
rect 94 -82 96 -80
rect 102 -82 104 -80
rect 122 -82 124 -80
rect 10 -98 12 -90
rect 10 -132 12 -102
rect 28 -110 30 -90
rect 36 -105 38 -90
rect 10 -137 12 -135
rect 28 -132 30 -114
rect 36 -132 38 -110
rect 52 -117 54 -90
rect 28 -137 30 -135
rect 36 -137 38 -135
rect 52 -132 54 -122
rect 69 -123 71 -90
rect 86 -104 88 -90
rect 52 -137 54 -135
rect 69 -132 71 -127
rect 69 -137 71 -135
rect 86 -132 88 -109
rect 94 -111 96 -90
rect 102 -106 104 -90
rect 122 -97 124 -90
rect 102 -109 107 -106
rect 91 -132 93 -116
rect 102 -119 104 -109
rect 96 -121 104 -119
rect 96 -132 98 -121
rect 86 -137 88 -135
rect 91 -137 93 -135
rect 96 -137 98 -135
rect 122 -132 124 -101
rect 122 -137 124 -135
<< polycontact >>
rect 26 107 30 111
rect 67 119 71 123
rect 50 113 54 118
rect 8 96 12 100
rect 35 102 39 107
rect 91 108 96 113
rect 84 101 88 106
rect 107 102 111 107
rect 120 94 124 98
rect 45 44 50 48
rect 56 33 60 38
rect 73 26 77 31
rect 98 50 103 54
rect 80 22 84 27
rect 108 40 113 44
rect 113 30 118 34
rect 118 14 123 18
rect 47 -31 51 -26
rect 45 -51 50 -47
rect 80 -36 84 -31
rect 73 -41 77 -36
rect 56 -48 60 -43
rect 8 -102 12 -98
rect 35 -110 39 -105
rect 26 -114 30 -110
rect 50 -122 54 -117
rect 84 -109 88 -104
rect 67 -127 71 -123
rect 91 -116 96 -111
rect 120 -101 124 -97
rect 107 -110 111 -105
<< metal1 >>
rect -2 144 157 146
rect -2 139 0 144
rect 5 139 9 144
rect 14 139 18 144
rect 23 139 27 144
rect 32 139 36 144
rect 41 139 45 144
rect 50 139 54 144
rect 59 139 63 144
rect 68 139 72 144
rect 77 139 81 144
rect 86 139 90 144
rect 95 139 99 144
rect 104 139 108 144
rect 113 139 117 144
rect 122 139 126 144
rect 131 139 135 144
rect 140 142 157 144
rect 140 139 149 142
rect -2 137 149 139
rect 154 137 157 142
rect 5 132 8 137
rect 23 132 26 137
rect 47 132 50 137
rect 64 132 67 137
rect 81 132 84 137
rect 117 132 120 137
rect 147 133 157 137
rect 15 111 18 127
rect 40 117 43 127
rect 57 123 60 127
rect 57 120 67 123
rect 40 114 50 117
rect 15 108 26 111
rect -1 96 8 99
rect 15 87 18 108
rect 43 99 46 114
rect 32 96 46 99
rect 32 87 35 96
rect 57 87 60 120
rect 74 113 77 127
rect 74 109 91 113
rect 74 87 77 109
rect 100 97 103 127
rect 127 102 130 127
rect 147 128 149 133
rect 154 128 157 133
rect 147 123 157 128
rect 147 118 149 123
rect 154 118 157 123
rect 147 113 157 118
rect 147 108 149 113
rect 154 108 157 113
rect 127 98 134 102
rect 147 101 157 108
rect 94 94 120 97
rect 90 87 93 93
rect 106 87 109 94
rect 127 87 130 98
rect 5 75 8 79
rect 23 75 26 79
rect 40 75 43 79
rect 147 96 149 101
rect 154 96 157 101
rect 147 89 157 96
rect 147 84 149 89
rect 154 84 157 89
rect 147 80 157 84
rect 47 75 50 79
rect 64 75 67 79
rect 82 75 85 79
rect 98 75 101 79
rect 117 75 120 79
rect 147 75 149 80
rect 154 75 157 80
rect -2 70 38 75
rect 43 70 47 75
rect 52 70 56 75
rect 61 70 65 75
rect 70 70 74 75
rect 79 70 83 75
rect 88 70 92 75
rect 97 70 101 75
rect 106 70 110 75
rect 115 70 119 75
rect 124 70 128 75
rect 133 70 140 75
rect 147 70 157 75
rect -2 69 27 70
rect -2 64 1 69
rect 6 64 10 69
rect 15 64 19 69
rect 24 64 27 69
rect -2 60 27 64
rect -2 55 1 60
rect 6 55 10 60
rect 15 55 19 60
rect 24 55 27 60
rect 43 66 46 70
rect 59 66 62 70
rect 71 66 74 70
rect 86 66 89 70
rect 98 66 101 70
rect 114 66 117 70
rect 130 66 133 70
rect 147 65 149 70
rect 154 65 157 70
rect 147 59 157 65
rect -2 52 27 55
rect 52 54 55 58
rect -2 49 10 52
rect 52 51 64 54
rect -2 44 1 49
rect 6 44 10 49
rect -2 39 10 44
rect -2 34 1 39
rect 6 34 10 39
rect -2 30 10 34
rect 65 30 68 51
rect 106 51 109 58
rect 122 51 125 58
rect 106 48 125 51
rect -2 25 1 30
rect 6 25 10 30
rect -2 21 10 25
rect -2 16 1 21
rect 6 16 10 21
rect -2 12 10 16
rect -2 7 1 12
rect 6 7 10 12
rect 60 27 73 30
rect 60 9 63 27
rect 122 26 125 48
rect 84 25 125 26
rect 147 54 149 59
rect 154 54 157 59
rect 147 50 157 54
rect 147 45 149 50
rect 154 45 157 50
rect 147 41 157 45
rect 147 36 149 41
rect 154 36 157 41
rect 147 32 157 36
rect 147 27 149 32
rect 154 27 157 32
rect 84 23 131 25
rect 122 22 131 23
rect 128 9 131 22
rect 147 23 157 27
rect 147 18 149 23
rect 154 18 157 23
rect 147 14 157 18
rect 147 9 149 14
rect 154 9 157 14
rect -2 3 10 7
rect -2 -2 1 3
rect 6 -2 10 3
rect 125 5 128 8
rect 147 5 157 9
rect 43 -2 46 4
rect 70 -2 73 4
rect 98 -2 101 4
rect 147 0 149 5
rect 154 0 157 5
rect 147 -2 157 0
rect -2 -6 10 -2
rect -2 -11 1 -6
rect 6 -11 10 -6
rect -2 -15 10 -11
rect 37 -5 157 -2
rect 37 -10 40 -5
rect 45 -10 49 -5
rect 54 -10 58 -5
rect 63 -10 67 -5
rect 72 -10 76 -5
rect 81 -10 85 -5
rect 90 -10 94 -5
rect 99 -10 103 -5
rect 108 -10 113 -5
rect 118 -10 140 -5
rect 145 -6 157 -5
rect 145 -10 149 -6
rect 37 -11 149 -10
rect 154 -11 157 -6
rect 37 -13 157 -11
rect -2 -20 1 -15
rect 6 -20 10 -15
rect -2 -25 10 -20
rect 43 -18 46 -13
rect 70 -18 73 -13
rect 147 -18 157 -13
rect 147 -23 148 -18
rect 153 -23 157 -18
rect -2 -30 1 -25
rect 6 -30 10 -25
rect -2 -35 10 -30
rect -2 -40 1 -35
rect 6 -40 10 -35
rect 60 -37 63 -23
rect 147 -30 157 -23
rect 84 -35 106 -32
rect 147 -35 148 -30
rect 153 -35 157 -30
rect 60 -40 73 -37
rect -2 -48 10 -40
rect -2 -53 1 -48
rect 6 -53 10 -48
rect 65 -52 68 -40
rect 147 -41 157 -35
rect -2 -55 10 -53
rect -2 -58 26 -55
rect -2 -63 1 -58
rect 6 -63 10 -58
rect 15 -63 19 -58
rect 24 -63 26 -58
rect 52 -57 64 -54
rect 147 -46 148 -41
rect 153 -46 157 -41
rect 147 -52 157 -46
rect 52 -61 55 -57
rect -2 -69 26 -63
rect -2 -74 1 -69
rect 6 -74 10 -69
rect 15 -74 19 -69
rect 24 -73 26 -69
rect 43 -73 46 -69
rect 59 -73 62 -69
rect 71 -73 74 -69
rect 87 -73 90 -69
rect 117 -64 140 -55
rect 117 -69 119 -64
rect 124 -69 128 -64
rect 133 -69 140 -64
rect 117 -73 140 -69
rect 24 -74 28 -73
rect -2 -78 28 -74
rect 33 -78 38 -73
rect 43 -78 47 -73
rect 52 -78 56 -73
rect 61 -78 65 -73
rect 70 -78 74 -73
rect 79 -78 83 -73
rect 88 -78 92 -73
rect 97 -78 101 -73
rect 106 -78 110 -73
rect 115 -78 119 -73
rect 124 -78 128 -73
rect 133 -78 140 -73
rect 147 -57 148 -52
rect 153 -57 157 -52
rect 147 -63 157 -57
rect 147 -68 148 -63
rect 153 -68 157 -63
rect 147 -73 157 -68
rect 147 -78 148 -73
rect 153 -78 157 -73
rect 5 -82 8 -78
rect 23 -82 26 -78
rect 40 -82 43 -78
rect 47 -82 50 -78
rect 64 -82 67 -78
rect 82 -82 85 -78
rect 98 -82 101 -78
rect 117 -82 120 -78
rect 0 -102 8 -99
rect 15 -111 18 -90
rect 32 -99 35 -90
rect 32 -102 46 -99
rect 15 -114 26 -111
rect 15 -131 18 -114
rect 43 -118 46 -102
rect 40 -121 50 -118
rect 40 -131 43 -121
rect 57 -124 60 -90
rect 74 -112 77 -90
rect 90 -96 93 -90
rect 106 -97 109 -90
rect 94 -100 120 -97
rect 74 -116 91 -112
rect 57 -127 67 -124
rect 57 -131 60 -127
rect 74 -131 77 -116
rect 100 -131 103 -100
rect 127 -101 130 -90
rect 147 -84 157 -78
rect 147 -89 148 -84
rect 153 -89 157 -84
rect 147 -94 157 -89
rect 147 -99 148 -94
rect 153 -99 157 -94
rect 127 -105 134 -101
rect 147 -104 157 -99
rect 127 -131 130 -105
rect 147 -109 148 -104
rect 153 -109 157 -104
rect 147 -114 157 -109
rect 147 -119 148 -114
rect 153 -119 157 -114
rect 147 -123 157 -119
rect 147 -128 148 -123
rect 153 -128 157 -123
rect 147 -132 157 -128
rect 5 -141 8 -136
rect 23 -141 26 -136
rect 47 -141 50 -136
rect 64 -141 67 -136
rect 81 -141 84 -136
rect 117 -141 120 -136
rect 147 -137 148 -132
rect 153 -137 157 -132
rect 147 -141 157 -137
rect -2 -143 157 -141
rect -2 -148 0 -143
rect 5 -148 9 -143
rect 14 -148 18 -143
rect 23 -148 27 -143
rect 32 -148 36 -143
rect 41 -148 45 -143
rect 50 -148 54 -143
rect 59 -148 63 -143
rect 68 -148 72 -143
rect 77 -148 81 -143
rect 86 -148 90 -143
rect 95 -148 99 -143
rect 104 -148 108 -143
rect 113 -148 117 -143
rect 122 -148 126 -143
rect 131 -148 135 -143
rect 140 -148 148 -143
rect 153 -148 157 -143
rect -2 -150 157 -148
<< m2contact >>
rect 35 102 39 107
rect 84 101 88 106
rect 89 93 94 98
rect 107 102 111 107
rect 31 79 35 87
rect 78 58 82 66
rect 106 58 110 66
rect 64 51 69 55
rect 45 44 50 48
rect 56 33 60 38
rect 98 50 103 54
rect 108 40 113 44
rect 118 14 123 18
rect 86 4 90 9
rect 128 4 133 9
rect 86 -23 90 -18
rect 47 -31 51 -26
rect 106 -36 110 -31
rect 45 -51 50 -47
rect 56 -48 60 -43
rect 64 -57 68 -52
rect 78 -69 82 -61
rect 31 -90 35 -82
rect 35 -110 39 -105
rect 89 -101 94 -96
rect 84 -109 88 -104
rect 107 -110 111 -105
<< metal2 >>
rect 39 103 67 106
rect 64 97 67 103
rect 64 94 89 97
rect 78 37 81 58
rect 60 34 90 37
rect 87 9 90 34
rect 87 -44 90 -23
rect 60 -47 90 -44
rect 78 -61 81 -47
rect 64 -100 89 -97
rect 64 -106 67 -100
rect 39 -109 67 -106
<< m3contact >>
rect 84 101 88 106
rect 107 102 111 107
rect 31 79 35 87
rect 106 58 110 66
rect 64 51 69 55
rect 45 44 50 48
rect 98 50 103 54
rect 108 40 113 44
rect 118 14 123 18
rect 128 4 133 9
rect 47 -31 51 -26
rect 45 -51 50 -47
rect 106 -36 110 -31
rect 64 -57 68 -52
rect 31 -90 35 -82
rect 84 -109 88 -104
rect 107 -110 111 -105
<< metal3 >>
rect 50 45 95 48
rect 92 43 95 45
rect 92 40 108 43
<< m4contact >>
rect 84 101 88 106
rect 107 102 111 107
rect 31 79 35 87
rect 106 58 110 66
rect 64 51 69 55
rect 98 50 103 54
rect 45 44 50 48
rect 118 14 123 18
rect 128 4 133 9
rect 47 -31 51 -26
rect 106 -36 110 -31
rect 45 -51 50 -47
rect 64 -57 68 -52
rect 31 -90 35 -82
rect 84 -109 88 -104
rect 107 -110 111 -105
<< metal4 >>
rect 78 102 84 105
rect 32 48 35 79
rect 78 74 81 102
rect 65 71 81 74
rect 65 55 68 71
rect 107 66 110 102
rect 69 51 98 54
rect 32 45 45 48
rect 93 14 118 17
rect 93 -27 96 14
rect 128 -20 131 4
rect 51 -30 96 -27
rect 107 -23 131 -20
rect 107 -31 110 -23
rect 32 -51 45 -48
rect 32 -82 35 -51
rect 65 -74 68 -57
rect 65 -77 81 -74
rect 78 -105 81 -77
rect 78 -108 84 -105
rect 107 -105 110 -36
<< labels >>
rlabel metal1 25 -147 25 -147 1 gnd!
rlabel metal1 134 -105 134 -101 1 dn
rlabel metal1 134 98 134 102 1 up
rlabel metal1 7 61 7 61 1 vdd!
rlabel metal1 -1 96 -1 99 3 fin
rlabel metal1 0 -102 0 -99 3 fvco_8
<< end >>
