magic
tech scmos
timestamp 1598983265
<< nwell >>
rect 0 0 146 25
<< ntransistor >>
rect 11 53 13 56
rect 28 53 30 56
rect 33 53 35 56
rect 49 53 51 56
rect 54 53 56 56
rect 70 53 72 56
rect 75 53 77 56
rect 91 53 93 56
rect 96 53 98 56
rect 112 53 114 56
rect 117 53 119 56
rect 133 53 135 56
<< ptransistor >>
rect 11 13 13 19
rect 28 13 30 19
rect 33 13 35 19
rect 49 13 51 19
rect 54 13 56 19
rect 70 13 72 19
rect 75 13 77 19
rect 91 13 93 19
rect 96 13 98 19
rect 112 13 114 19
rect 117 13 119 19
rect 133 13 135 19
<< ndiffusion >>
rect 10 53 11 56
rect 13 53 15 56
rect 27 53 28 56
rect 30 53 33 56
rect 35 53 36 56
rect 48 53 49 56
rect 51 53 54 56
rect 56 53 57 56
rect 69 53 70 56
rect 72 53 75 56
rect 77 53 78 56
rect 90 53 91 56
rect 93 53 96 56
rect 98 53 99 56
rect 111 53 112 56
rect 114 53 117 56
rect 119 53 120 56
rect 132 53 133 56
rect 135 53 136 56
<< pdiffusion >>
rect 10 13 11 19
rect 13 13 14 19
rect 27 13 28 19
rect 30 13 33 19
rect 35 13 36 19
rect 48 13 49 19
rect 51 13 54 19
rect 56 13 57 19
rect 69 13 70 19
rect 72 13 75 19
rect 77 13 78 19
rect 90 13 91 19
rect 93 13 96 19
rect 98 13 99 19
rect 111 13 112 19
rect 114 13 117 19
rect 119 13 120 19
rect 132 13 133 19
rect 135 13 136 19
<< ndcontact >>
rect 6 52 10 57
rect 15 52 19 57
rect 23 52 27 57
rect 36 52 40 57
rect 44 52 48 57
rect 57 52 61 57
rect 65 52 69 57
rect 78 52 82 57
rect 86 52 90 57
rect 99 52 103 57
rect 107 52 111 57
rect 120 52 124 57
rect 128 52 132 57
rect 136 52 140 57
<< pdcontact >>
rect 6 13 10 19
rect 14 13 18 19
rect 23 13 27 19
rect 36 13 40 19
rect 44 13 48 19
rect 57 13 61 19
rect 65 13 69 19
rect 78 13 82 19
rect 86 13 90 19
rect 99 13 103 19
rect 107 13 111 19
rect 120 13 124 19
rect 128 13 132 19
rect 136 13 140 19
<< psubstratepcontact >>
rect 0 61 4 66
rect 8 61 12 66
rect 16 61 20 66
rect 24 61 28 66
rect 32 61 36 66
rect 42 61 46 66
rect 50 61 54 66
rect 58 61 62 66
rect 73 61 77 66
rect 82 61 86 66
rect 91 61 95 66
rect 99 61 103 66
rect 107 61 111 66
rect 115 61 119 66
rect 124 61 128 66
rect 132 61 136 66
rect 142 61 146 66
<< nsubstratencontact >>
rect 3 3 7 8
rect 11 3 15 8
rect 19 3 23 8
rect 27 3 31 8
rect 35 3 39 8
rect 43 3 47 8
rect 51 3 55 8
rect 59 3 63 8
rect 67 3 71 8
rect 75 3 79 8
rect 83 3 87 8
rect 91 3 95 8
rect 99 3 103 8
rect 107 3 111 8
rect 115 3 119 8
rect 123 3 127 8
rect 131 3 135 8
rect 139 3 143 8
<< polysilicon >>
rect 11 56 13 58
rect 11 40 13 53
rect 28 56 30 58
rect 33 56 35 58
rect 28 41 30 53
rect 33 49 35 53
rect 49 56 51 58
rect 54 56 56 58
rect 33 44 34 49
rect 49 41 51 53
rect 54 49 56 53
rect 70 56 72 58
rect 75 56 77 58
rect 54 44 55 49
rect 70 41 72 53
rect 75 49 77 53
rect 91 56 93 58
rect 96 56 98 58
rect 75 44 76 49
rect 91 41 93 53
rect 96 49 98 53
rect 112 56 114 58
rect 117 56 119 58
rect 96 44 97 49
rect 11 35 12 40
rect 28 36 29 41
rect 49 36 50 41
rect 70 36 71 41
rect 91 36 92 41
rect 112 40 114 53
rect 117 49 119 53
rect 133 56 135 58
rect 133 49 135 53
rect 117 44 118 49
rect 133 44 134 49
rect 11 19 13 35
rect 28 19 30 36
rect 33 19 35 22
rect 49 19 51 36
rect 54 19 56 22
rect 70 19 72 36
rect 75 19 77 22
rect 91 19 93 36
rect 112 35 113 40
rect 96 19 98 22
rect 112 19 114 35
rect 117 19 119 22
rect 133 19 135 22
rect 11 11 13 13
rect 28 11 30 13
rect 33 11 35 13
rect 49 11 51 13
rect 54 11 56 13
rect 70 11 72 13
rect 75 11 77 13
rect 91 11 93 13
rect 96 11 98 13
rect 112 11 114 13
rect 117 11 119 13
rect 133 11 135 13
<< polycontact >>
rect 34 44 38 49
rect 55 44 59 49
rect 76 44 80 49
rect 97 44 101 49
rect 12 35 16 40
rect 29 36 33 41
rect 50 36 54 41
rect 71 36 75 41
rect 92 36 96 41
rect 118 44 122 49
rect 134 44 138 49
rect 33 22 37 27
rect 54 22 58 27
rect 75 22 79 27
rect 113 35 117 40
rect 96 22 100 27
rect 117 22 121 27
rect 131 22 135 27
<< metal1 >>
rect 4 61 8 66
rect 12 61 16 66
rect 20 61 24 66
rect 28 61 32 66
rect 36 61 42 66
rect 46 61 50 66
rect 54 61 58 66
rect 62 61 73 66
rect 77 61 82 66
rect 86 61 91 66
rect 95 61 99 66
rect 103 61 107 66
rect 111 61 115 66
rect 119 61 124 66
rect 128 61 132 66
rect 136 61 142 66
rect 16 57 19 61
rect 37 57 40 61
rect 58 57 61 61
rect 79 57 82 61
rect 100 57 103 61
rect 121 57 124 61
rect 137 57 140 61
rect 6 40 9 52
rect 23 40 26 52
rect 44 41 47 52
rect 65 41 68 52
rect 86 41 89 52
rect 107 41 110 52
rect 0 35 9 40
rect 16 35 22 40
rect 33 38 47 41
rect 6 19 9 35
rect 23 19 26 35
rect 44 19 47 38
rect 54 38 68 41
rect 65 19 68 38
rect 75 38 89 41
rect 86 19 89 38
rect 96 38 110 41
rect 107 19 110 38
rect 128 19 131 52
rect 138 44 146 49
rect 15 8 18 13
rect 37 8 40 13
rect 58 8 61 13
rect 79 8 82 13
rect 100 8 103 13
rect 121 8 124 13
rect 137 8 140 13
rect 0 3 3 8
rect 7 3 11 8
rect 15 3 19 8
rect 23 3 27 8
rect 31 3 35 8
rect 39 3 43 8
rect 47 3 51 8
rect 55 3 59 8
rect 63 3 67 8
rect 71 3 75 8
rect 79 3 83 8
rect 87 3 91 8
rect 95 3 99 8
rect 103 3 107 8
rect 111 3 115 8
rect 119 3 123 8
rect 127 3 131 8
rect 135 3 139 8
rect 143 3 146 8
rect 0 0 146 3
<< m2contact >>
rect 34 44 38 49
rect 55 44 59 49
rect 76 44 80 49
rect 97 44 101 49
rect 118 44 122 49
rect 22 35 26 40
rect 33 22 37 27
rect 54 22 58 27
rect 75 22 79 27
rect 96 22 100 27
rect 113 35 117 40
rect 117 22 121 27
rect 134 44 138 49
rect 131 22 135 27
<< metal2 >>
rect 38 44 55 49
rect 59 44 76 49
rect 80 44 97 49
rect 101 44 118 49
rect 122 44 134 49
rect 37 22 54 27
rect 58 22 75 27
rect 79 22 96 27
rect 100 22 117 27
rect 121 22 131 27
<< m3contact >>
rect 22 35 26 40
rect 113 35 117 40
<< m4contact >>
rect 22 35 26 40
rect 113 35 117 40
<< metal4 >>
rect 26 35 113 40
<< labels >>
rlabel metal1 0 35 0 40 3 fout
rlabel metal1 146 44 146 49 7 vin
rlabel metal1 73 2 73 2 1 vdd!
rlabel metal1 70 63 70 63 5 gnd!
<< end >>
