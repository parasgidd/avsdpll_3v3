magic
tech scmos
timestamp 1598444483
<< nwell >>
rect -4 -27 484 -2
<< ntransistor >>
rect 10 50 12 53
rect 29 50 31 53
rect 49 50 51 53
rect 61 50 63 53
rect 79 50 81 53
rect 95 50 97 53
rect 109 50 111 53
rect 122 50 124 53
rect 143 50 145 53
rect 173 50 175 53
rect 192 50 194 53
rect 212 50 214 53
rect 224 50 226 53
rect 242 50 244 53
rect 258 50 260 53
rect 272 50 274 53
rect 285 50 287 53
rect 306 50 308 53
rect 336 50 338 53
rect 355 50 357 53
rect 375 50 377 53
rect 387 50 389 53
rect 405 50 407 53
rect 421 50 423 53
rect 435 50 437 53
rect 448 50 450 53
rect 469 50 471 53
<< ptransistor >>
rect 10 -16 12 -8
rect 29 -16 31 -8
rect 49 -16 51 -8
rect 61 -16 63 -8
rect 79 -16 81 -8
rect 95 -16 97 -8
rect 109 -16 111 -8
rect 122 -16 124 -8
rect 143 -16 145 -8
rect 173 -16 175 -8
rect 192 -16 194 -8
rect 212 -16 214 -8
rect 224 -16 226 -8
rect 242 -16 244 -8
rect 258 -16 260 -8
rect 272 -16 274 -8
rect 285 -16 287 -8
rect 306 -16 308 -8
rect 336 -16 338 -8
rect 355 -16 357 -8
rect 375 -16 377 -8
rect 387 -16 389 -8
rect 405 -16 407 -8
rect 421 -16 423 -8
rect 435 -16 437 -8
rect 448 -16 450 -8
rect 469 -16 471 -8
<< ndiffusion >>
rect 7 50 10 53
rect 12 50 13 53
rect 27 50 29 53
rect 31 50 32 53
rect 46 50 49 53
rect 51 50 54 53
rect 59 50 61 53
rect 63 50 64 53
rect 78 50 79 53
rect 81 50 86 53
rect 91 50 95 53
rect 97 50 101 53
rect 106 50 109 53
rect 111 50 114 53
rect 119 50 122 53
rect 124 50 127 53
rect 141 50 143 53
rect 145 50 146 53
rect 170 50 173 53
rect 175 50 176 53
rect 190 50 192 53
rect 194 50 195 53
rect 209 50 212 53
rect 214 50 217 53
rect 222 50 224 53
rect 226 50 227 53
rect 241 50 242 53
rect 244 50 249 53
rect 254 50 258 53
rect 260 50 264 53
rect 269 50 272 53
rect 274 50 277 53
rect 282 50 285 53
rect 287 50 290 53
rect 304 50 306 53
rect 308 50 309 53
rect 333 50 336 53
rect 338 50 339 53
rect 353 50 355 53
rect 357 50 358 53
rect 372 50 375 53
rect 377 50 380 53
rect 385 50 387 53
rect 389 50 390 53
rect 404 50 405 53
rect 407 50 412 53
rect 417 50 421 53
rect 423 50 427 53
rect 432 50 435 53
rect 437 50 440 53
rect 445 50 448 53
rect 450 50 453 53
rect 467 50 469 53
rect 471 50 472 53
<< pdiffusion >>
rect 7 -16 10 -8
rect 12 -16 13 -8
rect 27 -16 29 -8
rect 31 -16 32 -8
rect 46 -16 49 -8
rect 51 -16 54 -8
rect 59 -16 61 -8
rect 63 -16 64 -8
rect 78 -16 79 -8
rect 81 -16 86 -8
rect 91 -16 95 -8
rect 97 -16 101 -8
rect 106 -16 109 -8
rect 111 -16 114 -8
rect 119 -16 122 -8
rect 124 -16 127 -8
rect 141 -16 143 -8
rect 145 -16 146 -8
rect 170 -16 173 -8
rect 175 -16 176 -8
rect 190 -16 192 -8
rect 194 -16 195 -8
rect 209 -16 212 -8
rect 214 -16 217 -8
rect 222 -16 224 -8
rect 226 -16 227 -8
rect 241 -16 242 -8
rect 244 -16 249 -8
rect 254 -16 258 -8
rect 260 -16 264 -8
rect 269 -16 272 -8
rect 274 -16 277 -8
rect 282 -16 285 -8
rect 287 -16 290 -8
rect 304 -16 306 -8
rect 308 -16 309 -8
rect 333 -16 336 -8
rect 338 -16 339 -8
rect 353 -16 355 -8
rect 357 -16 358 -8
rect 372 -16 375 -8
rect 377 -16 380 -8
rect 385 -16 387 -8
rect 389 -16 390 -8
rect 404 -16 405 -8
rect 407 -16 412 -8
rect 417 -16 421 -8
rect 423 -16 427 -8
rect 432 -16 435 -8
rect 437 -16 440 -8
rect 445 -16 448 -8
rect 450 -16 453 -8
rect 467 -16 469 -8
rect 471 -16 472 -8
<< ndcontact >>
rect 2 49 7 54
rect 13 49 18 54
rect 22 49 27 54
rect 32 49 37 54
rect 41 49 46 54
rect 54 49 59 54
rect 64 49 69 54
rect 73 49 78 54
rect 86 49 91 54
rect 101 49 106 54
rect 114 49 119 54
rect 127 49 132 54
rect 136 49 141 54
rect 146 49 151 54
rect 165 49 170 54
rect 176 49 181 54
rect 185 49 190 54
rect 195 49 200 54
rect 204 49 209 54
rect 217 49 222 54
rect 227 49 232 54
rect 236 49 241 54
rect 249 49 254 54
rect 264 49 269 54
rect 277 49 282 54
rect 290 49 295 54
rect 299 49 304 54
rect 309 49 314 54
rect 328 49 333 54
rect 339 49 344 54
rect 348 49 353 54
rect 358 49 363 54
rect 367 49 372 54
rect 380 49 385 54
rect 390 49 395 54
rect 399 49 404 54
rect 412 49 417 54
rect 427 49 432 54
rect 440 49 445 54
rect 453 49 458 54
rect 462 49 467 54
rect 472 49 477 54
<< pdcontact >>
rect 2 -16 7 -8
rect 13 -16 18 -8
rect 22 -16 27 -8
rect 32 -16 37 -8
rect 41 -16 46 -8
rect 54 -16 59 -8
rect 64 -16 69 -8
rect 73 -16 78 -8
rect 86 -16 91 -8
rect 101 -16 106 -8
rect 114 -16 119 -8
rect 127 -16 132 -8
rect 136 -16 141 -8
rect 146 -16 151 -8
rect 165 -16 170 -8
rect 176 -16 181 -8
rect 185 -16 190 -8
rect 195 -16 200 -8
rect 204 -16 209 -8
rect 217 -16 222 -8
rect 227 -16 232 -8
rect 236 -16 241 -8
rect 249 -16 254 -8
rect 264 -16 269 -8
rect 277 -16 282 -8
rect 290 -16 295 -8
rect 299 -16 304 -8
rect 309 -16 314 -8
rect 328 -16 333 -8
rect 339 -16 344 -8
rect 348 -16 353 -8
rect 358 -16 363 -8
rect 367 -16 372 -8
rect 380 -16 385 -8
rect 390 -16 395 -8
rect 399 -16 404 -8
rect 412 -16 417 -8
rect 427 -16 432 -8
rect 440 -16 445 -8
rect 453 -16 458 -8
rect 462 -16 467 -8
rect 472 -16 477 -8
<< psubstratepcontact >>
rect -2 80 3 85
rect 7 80 12 85
rect 16 80 21 85
rect 25 80 30 85
rect 35 80 40 85
rect 44 80 49 85
rect 54 80 59 85
rect 63 80 68 85
rect 74 80 79 85
rect 84 80 89 85
rect 93 80 98 85
rect 102 80 107 85
rect 111 80 116 85
rect 120 80 125 85
rect 129 80 134 85
rect 138 80 143 85
rect 147 80 152 85
rect 161 80 166 85
rect 170 80 175 85
rect 179 80 184 85
rect 188 80 193 85
rect 198 80 203 85
rect 207 80 212 85
rect 217 80 222 85
rect 226 80 231 85
rect 237 80 242 85
rect 247 80 252 85
rect 256 80 261 85
rect 265 80 270 85
rect 274 80 279 85
rect 283 80 288 85
rect 292 80 297 85
rect 301 80 306 85
rect 310 80 315 85
rect 324 80 329 85
rect 333 80 338 85
rect 342 80 347 85
rect 351 80 356 85
rect 361 80 366 85
rect 370 80 375 85
rect 380 80 385 85
rect 389 80 394 85
rect 400 80 405 85
rect 410 80 415 85
rect 419 80 424 85
rect 428 80 433 85
rect 437 80 442 85
rect 446 80 451 85
rect 455 80 460 85
rect 464 80 469 85
rect 473 80 478 85
rect -2 71 3 76
rect 7 71 12 76
rect 16 71 21 76
rect 25 71 30 76
rect 35 71 40 76
rect 44 71 49 76
rect 54 71 59 76
rect 63 71 68 76
rect 74 71 79 76
rect 84 71 89 76
rect 93 71 98 76
rect 102 71 107 76
rect 111 71 116 76
rect 120 71 125 76
rect 129 71 134 76
rect 138 71 143 76
rect 147 71 152 76
rect 161 71 166 76
rect 170 71 175 76
rect 179 71 184 76
rect 188 71 193 76
rect 198 71 203 76
rect 207 71 212 76
rect 217 71 222 76
rect 226 71 231 76
rect 237 71 242 76
rect 247 71 252 76
rect 256 71 261 76
rect 265 71 270 76
rect 274 71 279 76
rect 283 71 288 76
rect 292 71 297 76
rect 301 71 306 76
rect 310 71 315 76
rect 324 71 329 76
rect 333 71 338 76
rect 342 71 347 76
rect 351 71 356 76
rect 361 71 366 76
rect 370 71 375 76
rect 380 71 385 76
rect 389 71 394 76
rect 400 71 405 76
rect 410 71 415 76
rect 419 71 424 76
rect 428 71 433 76
rect 437 71 442 76
rect 446 71 451 76
rect 455 71 460 76
rect 464 71 469 76
rect 473 71 478 76
<< nsubstratencontact >>
rect -2 -42 3 -37
rect 7 -42 12 -37
rect 17 -42 22 -37
rect 26 -42 31 -37
rect 35 -42 40 -37
rect 44 -42 49 -37
rect 53 -42 58 -37
rect 62 -42 67 -37
rect 72 -42 77 -37
rect 81 -42 86 -37
rect 91 -42 96 -37
rect 101 -42 106 -37
rect 111 -42 116 -37
rect 120 -42 125 -37
rect 130 -42 135 -37
rect 139 -42 144 -37
rect 148 -42 153 -37
rect 161 -42 166 -37
rect 170 -42 175 -37
rect 180 -42 185 -37
rect 189 -42 194 -37
rect 198 -42 203 -37
rect 207 -42 212 -37
rect 216 -42 221 -37
rect 225 -42 230 -37
rect 235 -42 240 -37
rect 244 -42 249 -37
rect 254 -42 259 -37
rect 264 -42 269 -37
rect 274 -42 279 -37
rect 283 -42 288 -37
rect 293 -42 298 -37
rect 302 -42 307 -37
rect 311 -42 316 -37
rect 324 -42 329 -37
rect 333 -42 338 -37
rect 343 -42 348 -37
rect 352 -42 357 -37
rect 361 -42 366 -37
rect 370 -42 375 -37
rect 379 -42 384 -37
rect 388 -42 393 -37
rect 398 -42 403 -37
rect 407 -42 412 -37
rect 417 -42 422 -37
rect 427 -42 432 -37
rect 437 -42 442 -37
rect 446 -42 451 -37
rect 456 -42 461 -37
rect 465 -42 470 -37
rect 474 -42 479 -37
rect -2 -51 3 -46
rect 7 -51 12 -46
rect 17 -51 22 -46
rect 26 -51 31 -46
rect 35 -51 40 -46
rect 44 -51 49 -46
rect 53 -51 58 -46
rect 62 -51 67 -46
rect 72 -51 77 -46
rect 81 -51 86 -46
rect 91 -51 96 -46
rect 101 -51 106 -46
rect 111 -51 116 -46
rect 120 -51 125 -46
rect 130 -51 135 -46
rect 139 -51 144 -46
rect 148 -51 153 -46
rect 161 -51 166 -46
rect 170 -51 175 -46
rect 180 -51 185 -46
rect 189 -51 194 -46
rect 198 -51 203 -46
rect 207 -51 212 -46
rect 216 -51 221 -46
rect 225 -51 230 -46
rect 235 -51 240 -46
rect 244 -51 249 -46
rect 254 -51 259 -46
rect 264 -51 269 -46
rect 274 -51 279 -46
rect 283 -51 288 -46
rect 293 -51 298 -46
rect 302 -51 307 -46
rect 311 -51 316 -46
rect 324 -51 329 -46
rect 333 -51 338 -46
rect 343 -51 348 -46
rect 352 -51 357 -46
rect 361 -51 366 -46
rect 370 -51 375 -46
rect 379 -51 384 -46
rect 388 -51 393 -46
rect 398 -51 403 -46
rect 407 -51 412 -46
rect 417 -51 422 -46
rect 427 -51 432 -46
rect 437 -51 442 -46
rect 446 -51 451 -46
rect 456 -51 461 -46
rect 465 -51 470 -46
rect 474 -51 479 -46
<< polysilicon >>
rect 10 53 12 55
rect 10 7 12 50
rect 29 53 31 55
rect 29 17 31 50
rect 49 53 51 55
rect 49 32 51 50
rect 61 53 63 55
rect 10 -8 12 2
rect 29 -8 31 12
rect 61 10 63 50
rect 79 53 81 55
rect 79 48 81 50
rect 95 53 97 55
rect 95 48 97 50
rect 109 53 111 55
rect 79 46 97 48
rect 109 33 111 50
rect 122 53 124 55
rect 122 24 124 50
rect 143 53 145 55
rect 143 32 145 50
rect 173 53 175 55
rect 49 -8 51 -2
rect 61 -8 63 5
rect 79 -6 94 -4
rect 79 -8 81 -6
rect 95 -8 97 -6
rect 109 -8 111 -2
rect 122 -8 124 19
rect 143 -8 145 27
rect 173 7 175 50
rect 192 53 194 55
rect 192 17 194 50
rect 212 53 214 55
rect 212 32 214 50
rect 224 53 226 55
rect 173 -8 175 2
rect 192 -8 194 12
rect 224 10 226 50
rect 242 53 244 55
rect 242 48 244 50
rect 258 53 260 55
rect 258 48 260 50
rect 272 53 274 55
rect 242 46 260 48
rect 272 33 274 50
rect 285 53 287 55
rect 285 24 287 50
rect 306 53 308 55
rect 306 32 308 50
rect 336 53 338 55
rect 212 -8 214 -2
rect 224 -8 226 5
rect 242 -6 257 -4
rect 242 -8 244 -6
rect 258 -8 260 -6
rect 272 -8 274 -2
rect 285 -8 287 19
rect 306 -8 308 27
rect 336 7 338 50
rect 355 53 357 55
rect 355 17 357 50
rect 375 53 377 55
rect 375 32 377 50
rect 387 53 389 55
rect 336 -8 338 2
rect 355 -8 357 12
rect 387 10 389 50
rect 405 53 407 55
rect 405 48 407 50
rect 421 53 423 55
rect 421 48 423 50
rect 435 53 437 55
rect 405 46 423 48
rect 435 33 437 50
rect 448 53 450 55
rect 448 24 450 50
rect 469 53 471 55
rect 469 32 471 50
rect 375 -8 377 -2
rect 387 -8 389 5
rect 405 -6 420 -4
rect 405 -8 407 -6
rect 421 -8 423 -6
rect 435 -8 437 -2
rect 448 -8 450 19
rect 469 -8 471 27
rect 10 -18 12 -16
rect 29 -18 31 -16
rect 49 -18 51 -16
rect 61 -18 63 -16
rect 79 -18 81 -16
rect 95 -18 97 -16
rect 109 -18 111 -16
rect 122 -18 124 -16
rect 143 -18 145 -16
rect 173 -18 175 -16
rect 192 -18 194 -16
rect 212 -18 214 -16
rect 224 -18 226 -16
rect 242 -18 244 -16
rect 258 -18 260 -16
rect 272 -18 274 -16
rect 285 -18 287 -16
rect 306 -18 308 -16
rect 336 -18 338 -16
rect 355 -18 357 -16
rect 375 -18 377 -16
rect 387 -18 389 -16
rect 405 -18 407 -16
rect 421 -18 423 -16
rect 435 -18 437 -16
rect 448 -18 450 -16
rect 469 -18 471 -16
<< polycontact >>
rect 48 27 52 32
rect 29 12 33 17
rect 10 2 14 7
rect 80 41 84 46
rect 108 28 112 33
rect 143 27 147 32
rect 122 19 126 24
rect 61 5 65 10
rect 48 -2 52 3
rect 94 -6 98 -1
rect 108 -2 112 3
rect 211 27 215 32
rect 192 12 196 17
rect 173 2 177 7
rect 243 41 247 46
rect 271 28 275 33
rect 306 27 310 32
rect 285 19 289 24
rect 224 5 228 10
rect 211 -2 215 3
rect 257 -6 261 -1
rect 271 -2 275 3
rect 374 27 378 32
rect 355 12 359 17
rect 336 2 340 7
rect 406 41 410 46
rect 434 28 438 33
rect 469 27 473 32
rect 448 19 452 24
rect 387 5 391 10
rect 374 -2 378 3
rect 420 -6 424 -1
rect 434 -2 438 3
<< metal1 >>
rect -4 85 483 89
rect -4 80 -2 85
rect 3 80 7 85
rect 12 80 16 85
rect 21 80 25 85
rect 30 80 35 85
rect 40 80 44 85
rect 49 80 54 85
rect 59 80 63 85
rect 68 80 74 85
rect 79 80 84 85
rect 89 80 93 85
rect 98 80 102 85
rect 107 80 111 85
rect 116 80 120 85
rect 125 80 129 85
rect 134 80 138 85
rect 143 80 147 85
rect 152 80 161 85
rect 166 80 170 85
rect 175 80 179 85
rect 184 80 188 85
rect 193 80 198 85
rect 203 80 207 85
rect 212 80 217 85
rect 222 80 226 85
rect 231 80 237 85
rect 242 80 247 85
rect 252 80 256 85
rect 261 80 265 85
rect 270 80 274 85
rect 279 80 283 85
rect 288 80 292 85
rect 297 80 301 85
rect 306 80 310 85
rect 315 80 324 85
rect 329 80 333 85
rect 338 80 342 85
rect 347 80 351 85
rect 356 80 361 85
rect 366 80 370 85
rect 375 80 380 85
rect 385 80 389 85
rect 394 80 400 85
rect 405 80 410 85
rect 415 80 419 85
rect 424 80 428 85
rect 433 80 437 85
rect 442 80 446 85
rect 451 80 455 85
rect 460 80 464 85
rect 469 80 473 85
rect 478 80 483 85
rect -4 76 483 80
rect -4 71 -2 76
rect 3 71 7 76
rect 12 71 16 76
rect 21 71 25 76
rect 30 71 35 76
rect 40 71 44 76
rect 49 71 54 76
rect 59 71 63 76
rect 68 71 74 76
rect 79 71 84 76
rect 89 71 93 76
rect 98 71 102 76
rect 107 71 111 76
rect 116 71 120 76
rect 125 71 129 76
rect 134 71 138 76
rect 143 71 147 76
rect 152 71 161 76
rect 166 71 170 76
rect 175 71 179 76
rect 184 71 188 76
rect 193 71 198 76
rect 203 71 207 76
rect 212 71 217 76
rect 222 71 226 76
rect 231 71 237 76
rect 242 71 247 76
rect 252 71 256 76
rect 261 71 265 76
rect 270 71 274 76
rect 279 71 283 76
rect 288 71 292 76
rect 297 71 301 76
rect 306 71 310 76
rect 315 71 324 76
rect 329 71 333 76
rect 338 71 342 76
rect 347 71 351 76
rect 356 71 361 76
rect 366 71 370 76
rect 375 71 380 76
rect 385 71 389 76
rect 394 71 400 76
rect 405 71 410 76
rect 415 71 419 76
rect 424 71 428 76
rect 433 71 437 76
rect 442 71 446 76
rect 451 71 455 76
rect 460 71 464 76
rect 469 71 473 76
rect 478 71 483 76
rect -4 69 483 71
rect 14 54 17 69
rect 33 54 36 69
rect 65 54 68 69
rect 128 54 131 69
rect 147 54 150 69
rect 177 54 180 69
rect 196 54 199 69
rect 228 54 231 69
rect 291 54 294 69
rect 310 54 313 69
rect 340 54 343 69
rect 359 54 362 69
rect 391 54 394 69
rect 454 54 457 69
rect 473 54 476 69
rect 3 39 6 49
rect 3 -8 6 34
rect 23 7 26 49
rect 42 24 45 49
rect 14 3 22 6
rect 23 -8 26 2
rect 42 -8 45 19
rect 55 -8 58 49
rect 74 24 77 49
rect 87 38 90 49
rect 74 -8 77 19
rect 87 -8 90 33
rect 102 17 105 49
rect 102 -8 105 12
rect 115 10 118 49
rect 137 12 140 49
rect 166 39 169 49
rect 147 28 154 31
rect 115 -8 118 5
rect 137 -8 140 7
rect 166 -8 169 34
rect 186 7 189 49
rect 205 24 208 49
rect 177 3 185 6
rect 186 -8 189 2
rect 205 -8 208 19
rect 218 -8 221 49
rect 237 24 240 49
rect 250 38 253 49
rect 237 -8 240 19
rect 250 -8 253 33
rect 265 17 268 49
rect 265 -8 268 12
rect 278 10 281 49
rect 300 12 303 49
rect 329 39 332 49
rect 310 28 317 31
rect 278 -8 281 5
rect 300 -8 303 7
rect 329 -8 332 34
rect 349 7 352 49
rect 368 24 371 49
rect 340 3 348 6
rect 349 -8 352 2
rect 368 -8 371 19
rect 381 -8 384 49
rect 400 24 403 49
rect 413 38 416 49
rect 400 -8 403 19
rect 413 -8 416 33
rect 428 17 431 49
rect 428 -8 431 12
rect 441 10 444 49
rect 463 12 466 49
rect 473 28 477 31
rect 441 -8 444 5
rect 463 -8 466 7
rect 14 -35 17 -16
rect 33 -35 36 -16
rect 65 -35 68 -16
rect 128 -35 131 -16
rect 147 -35 150 -16
rect 177 -35 180 -16
rect 196 -35 199 -16
rect 228 -35 231 -16
rect 291 -35 294 -16
rect 310 -35 313 -16
rect 340 -35 343 -16
rect 359 -35 362 -16
rect 391 -35 394 -16
rect 454 -35 457 -16
rect 473 -35 476 -16
rect -4 -37 483 -35
rect -4 -42 -2 -37
rect 3 -42 7 -37
rect 12 -42 17 -37
rect 22 -42 26 -37
rect 31 -42 35 -37
rect 40 -42 44 -37
rect 49 -42 53 -37
rect 58 -42 62 -37
rect 67 -42 72 -37
rect 77 -42 81 -37
rect 86 -42 91 -37
rect 96 -42 101 -37
rect 106 -42 111 -37
rect 116 -42 120 -37
rect 125 -42 130 -37
rect 135 -42 139 -37
rect 144 -42 148 -37
rect 153 -42 161 -37
rect 166 -42 170 -37
rect 175 -42 180 -37
rect 185 -42 189 -37
rect 194 -42 198 -37
rect 203 -42 207 -37
rect 212 -42 216 -37
rect 221 -42 225 -37
rect 230 -42 235 -37
rect 240 -42 244 -37
rect 249 -42 254 -37
rect 259 -42 264 -37
rect 269 -42 274 -37
rect 279 -42 283 -37
rect 288 -42 293 -37
rect 298 -42 302 -37
rect 307 -42 311 -37
rect 316 -42 324 -37
rect 329 -42 333 -37
rect 338 -42 343 -37
rect 348 -42 352 -37
rect 357 -42 361 -37
rect 366 -42 370 -37
rect 375 -42 379 -37
rect 384 -42 388 -37
rect 393 -42 398 -37
rect 403 -42 407 -37
rect 412 -42 417 -37
rect 422 -42 427 -37
rect 432 -42 437 -37
rect 442 -42 446 -37
rect 451 -42 456 -37
rect 461 -42 465 -37
rect 470 -42 474 -37
rect 479 -42 483 -37
rect -4 -46 483 -42
rect -4 -51 -2 -46
rect 3 -51 7 -46
rect 12 -51 17 -46
rect 22 -51 26 -46
rect 31 -51 35 -46
rect 40 -51 44 -46
rect 49 -51 53 -46
rect 58 -51 62 -46
rect 67 -51 72 -46
rect 77 -51 81 -46
rect 86 -51 91 -46
rect 96 -51 101 -46
rect 106 -51 111 -46
rect 116 -51 120 -46
rect 125 -51 130 -46
rect 135 -51 139 -46
rect 144 -51 148 -46
rect 153 -51 161 -46
rect 166 -51 170 -46
rect 175 -51 180 -46
rect 185 -51 189 -46
rect 194 -51 198 -46
rect 203 -51 207 -46
rect 212 -51 216 -46
rect 221 -51 225 -46
rect 230 -51 235 -46
rect 240 -51 244 -46
rect 249 -51 254 -46
rect 259 -51 264 -46
rect 269 -51 274 -46
rect 279 -51 283 -46
rect 288 -51 293 -46
rect 298 -51 302 -46
rect 307 -51 311 -46
rect 316 -51 324 -46
rect 329 -51 333 -46
rect 338 -51 343 -46
rect 348 -51 352 -46
rect 357 -51 361 -46
rect 366 -51 370 -46
rect 375 -51 379 -46
rect 384 -51 388 -46
rect 393 -51 398 -46
rect 403 -51 407 -46
rect 412 -51 417 -46
rect 422 -51 427 -46
rect 432 -51 437 -46
rect 442 -51 446 -46
rect 451 -51 456 -46
rect 461 -51 465 -46
rect 470 -51 474 -46
rect 479 -51 483 -46
rect -4 -53 483 -51
<< m2contact >>
rect 3 34 7 39
rect 48 27 52 32
rect 42 19 46 24
rect 29 12 33 17
rect 10 2 14 7
rect 22 2 26 7
rect 48 -2 52 3
rect 80 41 84 46
rect 86 33 90 38
rect 73 19 77 24
rect 61 5 65 10
rect 108 28 112 33
rect 101 12 105 17
rect 94 -6 98 -1
rect 122 19 126 24
rect 166 34 170 39
rect 143 27 147 32
rect 154 26 158 31
rect 115 5 119 10
rect 136 7 140 12
rect 108 -2 112 3
rect 211 27 215 32
rect 205 19 209 24
rect 192 12 196 17
rect 173 2 177 7
rect 185 2 189 7
rect 211 -2 215 3
rect 243 41 247 46
rect 249 33 253 38
rect 236 19 240 24
rect 224 5 228 10
rect 271 28 275 33
rect 264 12 268 17
rect 257 -6 261 -1
rect 285 19 289 24
rect 329 34 333 39
rect 306 27 310 32
rect 317 26 321 31
rect 278 5 282 10
rect 299 7 303 12
rect 271 -2 275 3
rect 374 27 378 32
rect 368 19 372 24
rect 355 12 359 17
rect 336 2 340 7
rect 348 2 352 7
rect 374 -2 378 3
rect 406 41 410 46
rect 412 33 416 38
rect 399 19 403 24
rect 387 5 391 10
rect 434 28 438 33
rect 427 12 431 17
rect 420 -6 424 -1
rect 448 19 452 24
rect 469 27 473 32
rect 441 5 445 10
rect 462 7 466 12
rect 434 -2 438 3
<< metal2 >>
rect 7 35 86 38
rect 170 35 249 38
rect 333 35 412 38
rect 46 19 73 22
rect 77 20 122 23
rect 33 13 101 16
rect -6 3 10 6
rect 65 6 115 9
rect 155 6 158 26
rect 209 19 236 22
rect 240 20 285 23
rect 196 13 264 16
rect 155 3 173 6
rect 228 6 278 9
rect 318 6 321 26
rect 372 19 399 22
rect 403 20 448 23
rect 359 13 427 16
rect 318 3 336 6
rect 391 6 441 9
<< m3contact >>
rect 80 41 84 46
rect 243 41 247 46
rect 406 41 410 46
rect 48 27 52 32
rect 108 28 112 33
rect 143 27 147 32
rect 211 27 215 32
rect 271 28 275 33
rect 306 27 310 32
rect 374 27 378 32
rect 434 28 438 33
rect 469 27 473 32
rect 136 7 140 12
rect 48 -2 52 3
rect 94 -6 98 -1
rect 108 -2 112 3
rect 299 7 303 12
rect 211 -2 215 3
rect 257 -6 261 -1
rect 271 -2 275 3
rect 462 7 466 12
rect 374 -2 378 3
rect 420 -6 424 -1
rect 434 -2 438 3
<< metal3 >>
rect 52 28 108 31
rect 112 28 143 31
rect 94 -1 97 28
rect 215 28 271 31
rect 275 28 306 31
rect 257 -1 260 28
rect 378 28 434 31
rect 438 28 469 31
rect 420 -1 423 28
<< m4contact >>
rect 80 41 84 46
rect 243 41 247 46
rect 406 41 410 46
rect 48 -2 52 3
rect 136 7 140 12
rect 108 -2 112 3
rect 211 -2 215 3
rect 299 7 303 12
rect 271 -2 275 3
rect 374 -2 378 3
rect 462 7 466 12
rect 434 -2 438 3
<< metal4 >>
rect 80 11 83 41
rect 80 8 136 11
rect 80 3 83 8
rect 52 0 83 3
rect 108 3 111 8
rect 243 11 246 41
rect 243 8 299 11
rect 243 3 246 8
rect 215 0 246 3
rect 271 3 274 8
rect 406 11 409 41
rect 406 8 462 11
rect 406 3 409 8
rect 378 0 409 3
rect 434 3 437 8
<< labels >>
rlabel metal1 71 78 71 78 1 gnd!
rlabel metal2 -6 3 -6 6 3 q
rlabel metal1 234 78 234 78 1 gnd!
rlabel metal1 477 28 477 31 1 clk
rlabel metal1 397 78 397 78 1 gnd!
rlabel metal1 396 -45 396 -45 1 vdd!
rlabel metal1 233 -45 233 -45 1 vdd!
rlabel metal1 70 -45 70 -45 1 vdd!
<< end >>
