*__________________PLL-combined in 1 file_________________________*


XX1 f_in f_VCO/8 up down pfd_501
XX2 up down Vin_vco charge_pump
XX3 Vin_vco f_out vco_19_16
XX5 f_out N003 freq_div_2
XX6 N003 N002 freq_div_2
XX7 N002 f_VCO/8 freq_div_2
V1 f_in 0 PULSE 0 1.8 10p 60p 60p 100n 200n

.include osu018.lib

*V2 f_in 0 PULSE 0 1.8 10p 60p 60p 50n 100n
*V3 f_in 0 PULSE 0 1.8 10p 60p 60p 41.665n 83.33n

*___________LPF________________*
C1 Vin_vco 0 200p
C2 N001 0 500p
R1 Vin_vco N001 500
*______________________________*

*__________________Subcircuits_____________________*

******************PFD*******************************
.subckt pfd_501 f_clk_in f_VCO up down
XX1 N001 N005 N002 vddd 0 nand101
XX2 N002 N008 N006 vddd 0 nand101
XX3 N006 N007 N008 vddd 0 nand101
XX4 N007 N010 N011 vddd 0 nand101
XX5 N011 N009 N010 vddd 0 nand101
XX6 N013 N012 N009 vddd 0 nand101
XX7 f_clk_in N005 vddd 0 inv101
XX8 f_VCO N013 vddd 0 inv101
XX9 N002 N003 vddd 0 inv101
XX10 N003 N004 vddd 0 inv101
XX11 N009 N014 vddd 0 inv101
XX12 N014 N015 vddd 0 inv101
XX13 N004 N006 N007 N001 vddd 0 nand301
XX14 N007 N010 N015 N012 vddd 0 nand301
XX15 N012 down vddd 0 inv101
XX16 N006 N002 N009 N010 vddd 0 N007 nand401
XX17 N001 up vddd 0 inv101
V3 vddd 0 1.8
.ends pfd_501

*****************charge_pump*******************************
.subckt charge_pump UP Down CP
M7 UP_bar UP 0 0 nfet l=180n w=180n
M8 DOWN_bar Down 0 0 nfet l=180n w=180n
M12 VDD Down DOWN_bar VDD pfet l=180n w=540n
M14 VDD UP UP_bar VDD pfet l=180n w=540n
M15 UP_bar 0 N001 N001 nfet l=180n w=180n
M16 DOWN_bar 0 N004 N004 nfet l=180n w=180n
M17 N003 N004 N003 N003 nfet l=180n w=180n
M18 0 VDD VDD 0 nfet l=180n w=180n
M19 CP VDD N003 N003 nfet l=180n w=180n
M20 N003 Down 0 0 nfet l=180n w=15u
M21 N001 VDD UP_bar N001 pfet l=180n w=540n
M22 N004 VDD DOWN_bar N004 pfet l=180n w=540n
M23 N002 UP N002 N002 pfet l=180n w=540n
M24 0 0 VDD VDD pfet l=180n w=540n
M25 N002 0 CP N002 pfet l=180n w=540n
M26 VDD N001 N002 VDD pfet l=180n w=45u
V1 VDD 0 1.8
.ends charge_pump

******************VCO*******************************
.subckt vco_19_16 Vinvco osc
M7 Vp Vn 0 0 nfet l=180n w=360n
M8 Vp Vp VDD VDD pfet l=180n w=1800n
R1 Vn Vinvco 1
XU22 osc_fb Osc inv_20_10
XX3 n1 osc_fb Vp Vn cs_inv
XX16 N005 n1 Vp Vn cs_inv
XX17 N004 N005 Vp Vn cs_inv
XX18 N003 N004 Vp Vn cs_inv
XX19 N002 N003 Vp Vn cs_inv
XX20 N001 N002 Vp Vn cs_inv
XX21 osc_fb N001 Vp Vn cs_inv
V1 VDD 0 1.8
.ends vco_19_16

******************Frequency divider*******************************
.subckt freq_div_2 clock Q
M1 N004 N002 0 0 nfet l=180n w=180n
VDD VDD 0 1.8
M2 VDD N002 N004 VDD pfet l=180n w=540n
M5 N003 N004 0 0 nfet l=180n w=180n
M6 VDD N004 N003 VDD pfet l=180n w=540n
M7 D clock_b N002 0 nfet l=180n w=180n
M3 N002 clock D VDD pfet l=180n w=540n
M4 N002 clock N003 0 nfet l=180n w=180n
M8 N003 clock_b N002 VDD pfet l=180n w=540n
M9 Q N001 0 0 nfet l=180n w=180n
M10 VDD N001 Q VDD pfet l=180n w=540n
M11 D Q 0 0 nfet l=180n w=180n
M12 VDD Q D VDD pfet l=180n w=540n
M13 N004 clock N001 0 nfet l=180n w=180n
M14 N001 clock_b N004 VDD pfet l=180n w=540n
M15 N001 clock_b D 0 nfet l=180n w=180n
M16 D clock N001 VDD pfet l=180n w=540n
M17 clock_b clock 0 0 nfet l=180n w=180n
M18 VDD clock clock_b VDD pfet l=180n w=540n
.ends freq_div_2

.subckt nand101 in1 in2 out VDD GND
M1 out in1 N001 N001 nfet l=180n w=180n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 GND GND nfet l=180n w=360n
.ends nand101

.subckt inv101 in out VDD GND
M1 out in GND GND nfet l=180n w=180n
M2 VDD in out VDD pfet l=180n w=360n
.ends inv101

.subckt nand301 in1 in2 in3 out VDD GND
M1 out in1 N001 N001 nfet l=180n w=540n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 N002 N002 nfet l=180n w=540n
M5 N002 in3 GND GND nfet l=180n w=540n
M6 VDD in3 out VDD pfet l=180n w=360n
.ends nand301

.subckt nand401 in1 in2 in3 in4 VDD GND out
M1 out in1 N001 N001 nfet l=180n w=720n
M2 VDD in2 out VDD pfet l=180n w=360n
M3 VDD in1 out VDD pfet l=180n w=360n
M4 N001 in2 N002 N002 nfet l=180n w=720n
M5 N002 in3 N003 N003 nfet l=180n w=720n
M6 VDD in3 out VDD pfet l=180n w=360n
M7 N003 in4 GND GND nfet l=180n w=720n
M8 VDD in4 out VDD pfet l=180n w=360n
.ends nand401

.subckt inv_20_10 In Out
M1 Out In 0 0 nfet l=180n w=360n
M2 Out In N001 N001 pfet l=180n w=720n
V1 N001 0 1.8
.ends inv_20_10

.subckt cs_inv In Out Vp Vn
M1 N003 Vn 0 0 nfet l=180n w=360n
M4 N002 Vp N001 VDD pfet l=180n w=720n
M3 Out In N002 VDD pfet l=180n w=720n
M2 Out In N003 0 nfet l=180n w=360n
C1 Out 0 1f
V1 N001 0 1.8
.ends cs_inv


************simulation commands**************

.tran .1ns 6u
.ic V(vin_vco) = 0
.control
run
plot V(f_in)+8 V(up)+6 V(down)+4 V(Vin_vco)+2 V(f_out)

*plot V(N002)
*plot V(Vin_vco)
*plot V(f_out)
.endc
.end
